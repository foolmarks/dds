-----------------------------------------------------------------
--  File        : dpROM16_v1_0.vhd
--  Version     : 1
--  Revision    : 0
--  Date        : 12.03.2017
--  Author      : Mark Harvey
--  Description : Synchronous dual-port rom initialised to quarter sine wave
------------------------------------------------------------------


library ieee ;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;



entity dpROM16_v1_0 is
 port (
   CLK        : in  std_logic;          
   ADDRESS_A  : in  std_logic_vector;
   DATAOUT_A  : out std_logic_vector;
   ADDRESS_B  : in  std_logic_vector;
   DATAOUT_B  : out std_logic_vector
);
end entity dpROM16_v1_0;


architecture arcdpROM of dpROM16_v1_0 is

   signal dataA : std_logic_vector((DATAOUT_A'length -1) downto 0);
   signal dataB : std_logic_vector((DATAOUT_B'length -1) downto 0);

   type romType is array(0 to (2**ADDRESS_A'length)-1) of std_logic_vector((DATAOUT_A'length -1) downto 0);
   

   signal rom : romType := (
x"0000",x"0003",x"0006",x"0009",x"000D",x"0010",x"0013",x"0016",x"0019",x"001C",x"001F",x"0023",x"0026",x"0029",x"002C",x"002F",
x"0032",x"0035",x"0039",x"003C",x"003F",x"0042",x"0045",x"0048",x"004B",x"004F",x"0052",x"0055",x"0058",x"005B",x"005E",x"0061",
x"0065",x"0068",x"006B",x"006E",x"0071",x"0074",x"0077",x"007B",x"007E",x"0081",x"0084",x"0087",x"008A",x"008D",x"0091",x"0094",
x"0097",x"009A",x"009D",x"00A0",x"00A3",x"00A6",x"00AA",x"00AD",x"00B0",x"00B3",x"00B6",x"00B9",x"00BC",x"00C0",x"00C3",x"00C6",
x"00C9",x"00CC",x"00CF",x"00D2",x"00D6",x"00D9",x"00DC",x"00DF",x"00E2",x"00E5",x"00E8",x"00EC",x"00EF",x"00F2",x"00F5",x"00F8",
x"00FB",x"00FE",x"0102",x"0105",x"0108",x"010B",x"010E",x"0111",x"0114",x"0118",x"011B",x"011E",x"0121",x"0124",x"0127",x"012A",
x"012E",x"0131",x"0134",x"0137",x"013A",x"013D",x"0140",x"0144",x"0147",x"014A",x"014D",x"0150",x"0153",x"0156",x"015A",x"015D",
x"0160",x"0163",x"0166",x"0169",x"016C",x"0170",x"0173",x"0176",x"0179",x"017C",x"017F",x"0182",x"0186",x"0189",x"018C",x"018F",
x"0192",x"0195",x"0198",x"019C",x"019F",x"01A2",x"01A5",x"01A8",x"01AB",x"01AE",x"01B2",x"01B5",x"01B8",x"01BB",x"01BE",x"01C1",
x"01C4",x"01C8",x"01CB",x"01CE",x"01D1",x"01D4",x"01D7",x"01DA",x"01DD",x"01E1",x"01E4",x"01E7",x"01EA",x"01ED",x"01F0",x"01F3",
x"01F7",x"01FA",x"01FD",x"0200",x"0203",x"0206",x"0209",x"020D",x"0210",x"0213",x"0216",x"0219",x"021C",x"021F",x"0223",x"0226",
x"0229",x"022C",x"022F",x"0232",x"0235",x"0239",x"023C",x"023F",x"0242",x"0245",x"0248",x"024B",x"024F",x"0252",x"0255",x"0258",
x"025B",x"025E",x"0261",x"0265",x"0268",x"026B",x"026E",x"0271",x"0274",x"0277",x"027B",x"027E",x"0281",x"0284",x"0287",x"028A",
x"028D",x"0291",x"0294",x"0297",x"029A",x"029D",x"02A0",x"02A3",x"02A7",x"02AA",x"02AD",x"02B0",x"02B3",x"02B6",x"02B9",x"02BD",
x"02C0",x"02C3",x"02C6",x"02C9",x"02CC",x"02CF",x"02D2",x"02D6",x"02D9",x"02DC",x"02DF",x"02E2",x"02E5",x"02E8",x"02EC",x"02EF",
x"02F2",x"02F5",x"02F8",x"02FB",x"02FE",x"0302",x"0305",x"0308",x"030B",x"030E",x"0311",x"0314",x"0318",x"031B",x"031E",x"0321",
x"0324",x"0327",x"032A",x"032E",x"0331",x"0334",x"0337",x"033A",x"033D",x"0340",x"0344",x"0347",x"034A",x"034D",x"0350",x"0353",
x"0356",x"035A",x"035D",x"0360",x"0363",x"0366",x"0369",x"036C",x"0370",x"0373",x"0376",x"0379",x"037C",x"037F",x"0382",x"0385",
x"0389",x"038C",x"038F",x"0392",x"0395",x"0398",x"039B",x"039F",x"03A2",x"03A5",x"03A8",x"03AB",x"03AE",x"03B1",x"03B5",x"03B8",
x"03BB",x"03BE",x"03C1",x"03C4",x"03C7",x"03CB",x"03CE",x"03D1",x"03D4",x"03D7",x"03DA",x"03DD",x"03E1",x"03E4",x"03E7",x"03EA",
x"03ED",x"03F0",x"03F3",x"03F7",x"03FA",x"03FD",x"0400",x"0403",x"0406",x"0409",x"040D",x"0410",x"0413",x"0416",x"0419",x"041C",
x"041F",x"0423",x"0426",x"0429",x"042C",x"042F",x"0432",x"0435",x"0438",x"043C",x"043F",x"0442",x"0445",x"0448",x"044B",x"044E",
x"0452",x"0455",x"0458",x"045B",x"045E",x"0461",x"0464",x"0468",x"046B",x"046E",x"0471",x"0474",x"0477",x"047A",x"047E",x"0481",
x"0484",x"0487",x"048A",x"048D",x"0490",x"0494",x"0497",x"049A",x"049D",x"04A0",x"04A3",x"04A6",x"04AA",x"04AD",x"04B0",x"04B3",
x"04B6",x"04B9",x"04BC",x"04BF",x"04C3",x"04C6",x"04C9",x"04CC",x"04CF",x"04D2",x"04D5",x"04D9",x"04DC",x"04DF",x"04E2",x"04E5",
x"04E8",x"04EB",x"04EF",x"04F2",x"04F5",x"04F8",x"04FB",x"04FE",x"0501",x"0505",x"0508",x"050B",x"050E",x"0511",x"0514",x"0517",
x"051B",x"051E",x"0521",x"0524",x"0527",x"052A",x"052D",x"0530",x"0534",x"0537",x"053A",x"053D",x"0540",x"0543",x"0546",x"054A",
x"054D",x"0550",x"0553",x"0556",x"0559",x"055C",x"0560",x"0563",x"0566",x"0569",x"056C",x"056F",x"0572",x"0576",x"0579",x"057C",
x"057F",x"0582",x"0585",x"0588",x"058C",x"058F",x"0592",x"0595",x"0598",x"059B",x"059E",x"05A1",x"05A5",x"05A8",x"05AB",x"05AE",
x"05B1",x"05B4",x"05B7",x"05BB",x"05BE",x"05C1",x"05C4",x"05C7",x"05CA",x"05CD",x"05D1",x"05D4",x"05D7",x"05DA",x"05DD",x"05E0",
x"05E3",x"05E7",x"05EA",x"05ED",x"05F0",x"05F3",x"05F6",x"05F9",x"05FC",x"0600",x"0603",x"0606",x"0609",x"060C",x"060F",x"0612",
x"0616",x"0619",x"061C",x"061F",x"0622",x"0625",x"0628",x"062C",x"062F",x"0632",x"0635",x"0638",x"063B",x"063E",x"0642",x"0645",
x"0648",x"064B",x"064E",x"0651",x"0654",x"0657",x"065B",x"065E",x"0661",x"0664",x"0667",x"066A",x"066D",x"0671",x"0674",x"0677",
x"067A",x"067D",x"0680",x"0683",x"0687",x"068A",x"068D",x"0690",x"0693",x"0696",x"0699",x"069D",x"06A0",x"06A3",x"06A6",x"06A9",
x"06AC",x"06AF",x"06B2",x"06B6",x"06B9",x"06BC",x"06BF",x"06C2",x"06C5",x"06C8",x"06CC",x"06CF",x"06D2",x"06D5",x"06D8",x"06DB",
x"06DE",x"06E2",x"06E5",x"06E8",x"06EB",x"06EE",x"06F1",x"06F4",x"06F7",x"06FB",x"06FE",x"0701",x"0704",x"0707",x"070A",x"070D",
x"0711",x"0714",x"0717",x"071A",x"071D",x"0720",x"0723",x"0727",x"072A",x"072D",x"0730",x"0733",x"0736",x"0739",x"073C",x"0740",
x"0743",x"0746",x"0749",x"074C",x"074F",x"0752",x"0756",x"0759",x"075C",x"075F",x"0762",x"0765",x"0768",x"076C",x"076F",x"0772",
x"0775",x"0778",x"077B",x"077E",x"0781",x"0785",x"0788",x"078B",x"078E",x"0791",x"0794",x"0797",x"079B",x"079E",x"07A1",x"07A4",
x"07A7",x"07AA",x"07AD",x"07B1",x"07B4",x"07B7",x"07BA",x"07BD",x"07C0",x"07C3",x"07C6",x"07CA",x"07CD",x"07D0",x"07D3",x"07D6",
x"07D9",x"07DC",x"07E0",x"07E3",x"07E6",x"07E9",x"07EC",x"07EF",x"07F2",x"07F6",x"07F9",x"07FC",x"07FF",x"0802",x"0805",x"0808",
x"080B",x"080F",x"0812",x"0815",x"0818",x"081B",x"081E",x"0821",x"0825",x"0828",x"082B",x"082E",x"0831",x"0834",x"0837",x"083A",
x"083E",x"0841",x"0844",x"0847",x"084A",x"084D",x"0850",x"0854",x"0857",x"085A",x"085D",x"0860",x"0863",x"0866",x"086A",x"086D",
x"0870",x"0873",x"0876",x"0879",x"087C",x"087F",x"0883",x"0886",x"0889",x"088C",x"088F",x"0892",x"0895",x"0899",x"089C",x"089F",
x"08A2",x"08A5",x"08A8",x"08AB",x"08AE",x"08B2",x"08B5",x"08B8",x"08BB",x"08BE",x"08C1",x"08C4",x"08C8",x"08CB",x"08CE",x"08D1",
x"08D4",x"08D7",x"08DA",x"08DD",x"08E1",x"08E4",x"08E7",x"08EA",x"08ED",x"08F0",x"08F3",x"08F7",x"08FA",x"08FD",x"0900",x"0903",
x"0906",x"0909",x"090C",x"0910",x"0913",x"0916",x"0919",x"091C",x"091F",x"0922",x"0926",x"0929",x"092C",x"092F",x"0932",x"0935",
x"0938",x"093B",x"093F",x"0942",x"0945",x"0948",x"094B",x"094E",x"0951",x"0955",x"0958",x"095B",x"095E",x"0961",x"0964",x"0967",
x"096A",x"096E",x"0971",x"0974",x"0977",x"097A",x"097D",x"0980",x"0984",x"0987",x"098A",x"098D",x"0990",x"0993",x"0996",x"0999",
x"099D",x"09A0",x"09A3",x"09A6",x"09A9",x"09AC",x"09AF",x"09B3",x"09B6",x"09B9",x"09BC",x"09BF",x"09C2",x"09C5",x"09C8",x"09CC",
x"09CF",x"09D2",x"09D5",x"09D8",x"09DB",x"09DE",x"09E2",x"09E5",x"09E8",x"09EB",x"09EE",x"09F1",x"09F4",x"09F7",x"09FB",x"09FE",
x"0A01",x"0A04",x"0A07",x"0A0A",x"0A0D",x"0A11",x"0A14",x"0A17",x"0A1A",x"0A1D",x"0A20",x"0A23",x"0A26",x"0A2A",x"0A2D",x"0A30",
x"0A33",x"0A36",x"0A39",x"0A3C",x"0A3F",x"0A43",x"0A46",x"0A49",x"0A4C",x"0A4F",x"0A52",x"0A55",x"0A59",x"0A5C",x"0A5F",x"0A62",
x"0A65",x"0A68",x"0A6B",x"0A6E",x"0A72",x"0A75",x"0A78",x"0A7B",x"0A7E",x"0A81",x"0A84",x"0A87",x"0A8B",x"0A8E",x"0A91",x"0A94",
x"0A97",x"0A9A",x"0A9D",x"0AA1",x"0AA4",x"0AA7",x"0AAA",x"0AAD",x"0AB0",x"0AB3",x"0AB6",x"0ABA",x"0ABD",x"0AC0",x"0AC3",x"0AC6",
x"0AC9",x"0ACC",x"0ACF",x"0AD3",x"0AD6",x"0AD9",x"0ADC",x"0ADF",x"0AE2",x"0AE5",x"0AE9",x"0AEC",x"0AEF",x"0AF2",x"0AF5",x"0AF8",
x"0AFB",x"0AFE",x"0B02",x"0B05",x"0B08",x"0B0B",x"0B0E",x"0B11",x"0B14",x"0B17",x"0B1B",x"0B1E",x"0B21",x"0B24",x"0B27",x"0B2A",
x"0B2D",x"0B31",x"0B34",x"0B37",x"0B3A",x"0B3D",x"0B40",x"0B43",x"0B46",x"0B4A",x"0B4D",x"0B50",x"0B53",x"0B56",x"0B59",x"0B5C",
x"0B5F",x"0B63",x"0B66",x"0B69",x"0B6C",x"0B6F",x"0B72",x"0B75",x"0B78",x"0B7C",x"0B7F",x"0B82",x"0B85",x"0B88",x"0B8B",x"0B8E",
x"0B92",x"0B95",x"0B98",x"0B9B",x"0B9E",x"0BA1",x"0BA4",x"0BA7",x"0BAB",x"0BAE",x"0BB1",x"0BB4",x"0BB7",x"0BBA",x"0BBD",x"0BC0",
x"0BC4",x"0BC7",x"0BCA",x"0BCD",x"0BD0",x"0BD3",x"0BD6",x"0BD9",x"0BDD",x"0BE0",x"0BE3",x"0BE6",x"0BE9",x"0BEC",x"0BEF",x"0BF3",
x"0BF6",x"0BF9",x"0BFC",x"0BFF",x"0C02",x"0C05",x"0C08",x"0C0C",x"0C0F",x"0C12",x"0C15",x"0C18",x"0C1B",x"0C1E",x"0C21",x"0C25",
x"0C28",x"0C2B",x"0C2E",x"0C31",x"0C34",x"0C37",x"0C3A",x"0C3E",x"0C41",x"0C44",x"0C47",x"0C4A",x"0C4D",x"0C50",x"0C53",x"0C57",
x"0C5A",x"0C5D",x"0C60",x"0C63",x"0C66",x"0C69",x"0C6C",x"0C70",x"0C73",x"0C76",x"0C79",x"0C7C",x"0C7F",x"0C82",x"0C85",x"0C89",
x"0C8C",x"0C8F",x"0C92",x"0C95",x"0C98",x"0C9B",x"0C9E",x"0CA2",x"0CA5",x"0CA8",x"0CAB",x"0CAE",x"0CB1",x"0CB4",x"0CB7",x"0CBB",
x"0CBE",x"0CC1",x"0CC4",x"0CC7",x"0CCA",x"0CCD",x"0CD1",x"0CD4",x"0CD7",x"0CDA",x"0CDD",x"0CE0",x"0CE3",x"0CE6",x"0CEA",x"0CED",
x"0CF0",x"0CF3",x"0CF6",x"0CF9",x"0CFC",x"0CFF",x"0D03",x"0D06",x"0D09",x"0D0C",x"0D0F",x"0D12",x"0D15",x"0D18",x"0D1C",x"0D1F",
x"0D22",x"0D25",x"0D28",x"0D2B",x"0D2E",x"0D31",x"0D35",x"0D38",x"0D3B",x"0D3E",x"0D41",x"0D44",x"0D47",x"0D4A",x"0D4E",x"0D51",
x"0D54",x"0D57",x"0D5A",x"0D5D",x"0D60",x"0D63",x"0D66",x"0D6A",x"0D6D",x"0D70",x"0D73",x"0D76",x"0D79",x"0D7C",x"0D7F",x"0D83",
x"0D86",x"0D89",x"0D8C",x"0D8F",x"0D92",x"0D95",x"0D98",x"0D9C",x"0D9F",x"0DA2",x"0DA5",x"0DA8",x"0DAB",x"0DAE",x"0DB1",x"0DB5",
x"0DB8",x"0DBB",x"0DBE",x"0DC1",x"0DC4",x"0DC7",x"0DCA",x"0DCE",x"0DD1",x"0DD4",x"0DD7",x"0DDA",x"0DDD",x"0DE0",x"0DE3",x"0DE7",
x"0DEA",x"0DED",x"0DF0",x"0DF3",x"0DF6",x"0DF9",x"0DFC",x"0E00",x"0E03",x"0E06",x"0E09",x"0E0C",x"0E0F",x"0E12",x"0E15",x"0E19",
x"0E1C",x"0E1F",x"0E22",x"0E25",x"0E28",x"0E2B",x"0E2E",x"0E32",x"0E35",x"0E38",x"0E3B",x"0E3E",x"0E41",x"0E44",x"0E47",x"0E4A",
x"0E4E",x"0E51",x"0E54",x"0E57",x"0E5A",x"0E5D",x"0E60",x"0E63",x"0E67",x"0E6A",x"0E6D",x"0E70",x"0E73",x"0E76",x"0E79",x"0E7C",
x"0E80",x"0E83",x"0E86",x"0E89",x"0E8C",x"0E8F",x"0E92",x"0E95",x"0E99",x"0E9C",x"0E9F",x"0EA2",x"0EA5",x"0EA8",x"0EAB",x"0EAE",
x"0EB1",x"0EB5",x"0EB8",x"0EBB",x"0EBE",x"0EC1",x"0EC4",x"0EC7",x"0ECA",x"0ECE",x"0ED1",x"0ED4",x"0ED7",x"0EDA",x"0EDD",x"0EE0",
x"0EE3",x"0EE7",x"0EEA",x"0EED",x"0EF0",x"0EF3",x"0EF6",x"0EF9",x"0EFC",x"0EFF",x"0F03",x"0F06",x"0F09",x"0F0C",x"0F0F",x"0F12",
x"0F15",x"0F18",x"0F1C",x"0F1F",x"0F22",x"0F25",x"0F28",x"0F2B",x"0F2E",x"0F31",x"0F35",x"0F38",x"0F3B",x"0F3E",x"0F41",x"0F44",
x"0F47",x"0F4A",x"0F4D",x"0F51",x"0F54",x"0F57",x"0F5A",x"0F5D",x"0F60",x"0F63",x"0F66",x"0F6A",x"0F6D",x"0F70",x"0F73",x"0F76",
x"0F79",x"0F7C",x"0F7F",x"0F82",x"0F86",x"0F89",x"0F8C",x"0F8F",x"0F92",x"0F95",x"0F98",x"0F9B",x"0F9F",x"0FA2",x"0FA5",x"0FA8",
x"0FAB",x"0FAE",x"0FB1",x"0FB4",x"0FB8",x"0FBB",x"0FBE",x"0FC1",x"0FC4",x"0FC7",x"0FCA",x"0FCD",x"0FD0",x"0FD4",x"0FD7",x"0FDA",
x"0FDD",x"0FE0",x"0FE3",x"0FE6",x"0FE9",x"0FEC",x"0FF0",x"0FF3",x"0FF6",x"0FF9",x"0FFC",x"0FFF",x"1002",x"1005",x"1009",x"100C",
x"100F",x"1012",x"1015",x"1018",x"101B",x"101E",x"1021",x"1025",x"1028",x"102B",x"102E",x"1031",x"1034",x"1037",x"103A",x"103E",
x"1041",x"1044",x"1047",x"104A",x"104D",x"1050",x"1053",x"1056",x"105A",x"105D",x"1060",x"1063",x"1066",x"1069",x"106C",x"106F",
x"1072",x"1076",x"1079",x"107C",x"107F",x"1082",x"1085",x"1088",x"108B",x"108F",x"1092",x"1095",x"1098",x"109B",x"109E",x"10A1",
x"10A4",x"10A7",x"10AB",x"10AE",x"10B1",x"10B4",x"10B7",x"10BA",x"10BD",x"10C0",x"10C3",x"10C7",x"10CA",x"10CD",x"10D0",x"10D3",
x"10D6",x"10D9",x"10DC",x"10E0",x"10E3",x"10E6",x"10E9",x"10EC",x"10EF",x"10F2",x"10F5",x"10F8",x"10FC",x"10FF",x"1102",x"1105",
x"1108",x"110B",x"110E",x"1111",x"1114",x"1118",x"111B",x"111E",x"1121",x"1124",x"1127",x"112A",x"112D",x"1130",x"1134",x"1137",
x"113A",x"113D",x"1140",x"1143",x"1146",x"1149",x"114C",x"1150",x"1153",x"1156",x"1159",x"115C",x"115F",x"1162",x"1165",x"1168",
x"116C",x"116F",x"1172",x"1175",x"1178",x"117B",x"117E",x"1181",x"1185",x"1188",x"118B",x"118E",x"1191",x"1194",x"1197",x"119A",
x"119D",x"11A1",x"11A4",x"11A7",x"11AA",x"11AD",x"11B0",x"11B3",x"11B6",x"11B9",x"11BD",x"11C0",x"11C3",x"11C6",x"11C9",x"11CC",
x"11CF",x"11D2",x"11D5",x"11D9",x"11DC",x"11DF",x"11E2",x"11E5",x"11E8",x"11EB",x"11EE",x"11F1",x"11F5",x"11F8",x"11FB",x"11FE",
x"1201",x"1204",x"1207",x"120A",x"120D",x"1210",x"1214",x"1217",x"121A",x"121D",x"1220",x"1223",x"1226",x"1229",x"122C",x"1230",
x"1233",x"1236",x"1239",x"123C",x"123F",x"1242",x"1245",x"1248",x"124C",x"124F",x"1252",x"1255",x"1258",x"125B",x"125E",x"1261",
x"1264",x"1268",x"126B",x"126E",x"1271",x"1274",x"1277",x"127A",x"127D",x"1280",x"1284",x"1287",x"128A",x"128D",x"1290",x"1293",
x"1296",x"1299",x"129C",x"12A0",x"12A3",x"12A6",x"12A9",x"12AC",x"12AF",x"12B2",x"12B5",x"12B8",x"12BB",x"12BF",x"12C2",x"12C5",
x"12C8",x"12CB",x"12CE",x"12D1",x"12D4",x"12D7",x"12DB",x"12DE",x"12E1",x"12E4",x"12E7",x"12EA",x"12ED",x"12F0",x"12F3",x"12F7",
x"12FA",x"12FD",x"1300",x"1303",x"1306",x"1309",x"130C",x"130F",x"1312",x"1316",x"1319",x"131C",x"131F",x"1322",x"1325",x"1328",
x"132B",x"132E",x"1332",x"1335",x"1338",x"133B",x"133E",x"1341",x"1344",x"1347",x"134A",x"134D",x"1351",x"1354",x"1357",x"135A",
x"135D",x"1360",x"1363",x"1366",x"1369",x"136D",x"1370",x"1373",x"1376",x"1379",x"137C",x"137F",x"1382",x"1385",x"1388",x"138C",
x"138F",x"1392",x"1395",x"1398",x"139B",x"139E",x"13A1",x"13A4",x"13A8",x"13AB",x"13AE",x"13B1",x"13B4",x"13B7",x"13BA",x"13BD",
x"13C0",x"13C3",x"13C7",x"13CA",x"13CD",x"13D0",x"13D3",x"13D6",x"13D9",x"13DC",x"13DF",x"13E3",x"13E6",x"13E9",x"13EC",x"13EF",
x"13F2",x"13F5",x"13F8",x"13FB",x"13FE",x"1402",x"1405",x"1408",x"140B",x"140E",x"1411",x"1414",x"1417",x"141A",x"141D",x"1421",
x"1424",x"1427",x"142A",x"142D",x"1430",x"1433",x"1436",x"1439",x"143C",x"1440",x"1443",x"1446",x"1449",x"144C",x"144F",x"1452",
x"1455",x"1458",x"145C",x"145F",x"1462",x"1465",x"1468",x"146B",x"146E",x"1471",x"1474",x"1477",x"147B",x"147E",x"1481",x"1484",
x"1487",x"148A",x"148D",x"1490",x"1493",x"1496",x"149A",x"149D",x"14A0",x"14A3",x"14A6",x"14A9",x"14AC",x"14AF",x"14B2",x"14B5",
x"14B9",x"14BC",x"14BF",x"14C2",x"14C5",x"14C8",x"14CB",x"14CE",x"14D1",x"14D4",x"14D8",x"14DB",x"14DE",x"14E1",x"14E4",x"14E7",
x"14EA",x"14ED",x"14F0",x"14F3",x"14F7",x"14FA",x"14FD",x"1500",x"1503",x"1506",x"1509",x"150C",x"150F",x"1512",x"1516",x"1519",
x"151C",x"151F",x"1522",x"1525",x"1528",x"152B",x"152E",x"1531",x"1534",x"1538",x"153B",x"153E",x"1541",x"1544",x"1547",x"154A",
x"154D",x"1550",x"1553",x"1557",x"155A",x"155D",x"1560",x"1563",x"1566",x"1569",x"156C",x"156F",x"1572",x"1576",x"1579",x"157C",
x"157F",x"1582",x"1585",x"1588",x"158B",x"158E",x"1591",x"1595",x"1598",x"159B",x"159E",x"15A1",x"15A4",x"15A7",x"15AA",x"15AD",
x"15B0",x"15B3",x"15B7",x"15BA",x"15BD",x"15C0",x"15C3",x"15C6",x"15C9",x"15CC",x"15CF",x"15D2",x"15D6",x"15D9",x"15DC",x"15DF",
x"15E2",x"15E5",x"15E8",x"15EB",x"15EE",x"15F1",x"15F4",x"15F8",x"15FB",x"15FE",x"1601",x"1604",x"1607",x"160A",x"160D",x"1610",
x"1613",x"1617",x"161A",x"161D",x"1620",x"1623",x"1626",x"1629",x"162C",x"162F",x"1632",x"1635",x"1639",x"163C",x"163F",x"1642",
x"1645",x"1648",x"164B",x"164E",x"1651",x"1654",x"1657",x"165B",x"165E",x"1661",x"1664",x"1667",x"166A",x"166D",x"1670",x"1673",
x"1676",x"167A",x"167D",x"1680",x"1683",x"1686",x"1689",x"168C",x"168F",x"1692",x"1695",x"1698",x"169C",x"169F",x"16A2",x"16A5",
x"16A8",x"16AB",x"16AE",x"16B1",x"16B4",x"16B7",x"16BA",x"16BE",x"16C1",x"16C4",x"16C7",x"16CA",x"16CD",x"16D0",x"16D3",x"16D6",
x"16D9",x"16DC",x"16E0",x"16E3",x"16E6",x"16E9",x"16EC",x"16EF",x"16F2",x"16F5",x"16F8",x"16FB",x"16FE",x"1702",x"1705",x"1708",
x"170B",x"170E",x"1711",x"1714",x"1717",x"171A",x"171D",x"1720",x"1724",x"1727",x"172A",x"172D",x"1730",x"1733",x"1736",x"1739",
x"173C",x"173F",x"1742",x"1746",x"1749",x"174C",x"174F",x"1752",x"1755",x"1758",x"175B",x"175E",x"1761",x"1764",x"1767",x"176B",
x"176E",x"1771",x"1774",x"1777",x"177A",x"177D",x"1780",x"1783",x"1786",x"1789",x"178D",x"1790",x"1793",x"1796",x"1799",x"179C",
x"179F",x"17A2",x"17A5",x"17A8",x"17AB",x"17AF",x"17B2",x"17B5",x"17B8",x"17BB",x"17BE",x"17C1",x"17C4",x"17C7",x"17CA",x"17CD",
x"17D0",x"17D4",x"17D7",x"17DA",x"17DD",x"17E0",x"17E3",x"17E6",x"17E9",x"17EC",x"17EF",x"17F2",x"17F6",x"17F9",x"17FC",x"17FF",
x"1802",x"1805",x"1808",x"180B",x"180E",x"1811",x"1814",x"1817",x"181B",x"181E",x"1821",x"1824",x"1827",x"182A",x"182D",x"1830",
x"1833",x"1836",x"1839",x"183C",x"1840",x"1843",x"1846",x"1849",x"184C",x"184F",x"1852",x"1855",x"1858",x"185B",x"185E",x"1861",
x"1865",x"1868",x"186B",x"186E",x"1871",x"1874",x"1877",x"187A",x"187D",x"1880",x"1883",x"1886",x"188A",x"188D",x"1890",x"1893",
x"1896",x"1899",x"189C",x"189F",x"18A2",x"18A5",x"18A8",x"18AB",x"18AF",x"18B2",x"18B5",x"18B8",x"18BB",x"18BE",x"18C1",x"18C4",
x"18C7",x"18CA",x"18CD",x"18D0",x"18D4",x"18D7",x"18DA",x"18DD",x"18E0",x"18E3",x"18E6",x"18E9",x"18EC",x"18EF",x"18F2",x"18F5",
x"18F9",x"18FC",x"18FF",x"1902",x"1905",x"1908",x"190B",x"190E",x"1911",x"1914",x"1917",x"191A",x"191D",x"1921",x"1924",x"1927",
x"192A",x"192D",x"1930",x"1933",x"1936",x"1939",x"193C",x"193F",x"1942",x"1946",x"1949",x"194C",x"194F",x"1952",x"1955",x"1958",
x"195B",x"195E",x"1961",x"1964",x"1967",x"196A",x"196E",x"1971",x"1974",x"1977",x"197A",x"197D",x"1980",x"1983",x"1986",x"1989",
x"198C",x"198F",x"1993",x"1996",x"1999",x"199C",x"199F",x"19A2",x"19A5",x"19A8",x"19AB",x"19AE",x"19B1",x"19B4",x"19B7",x"19BB",
x"19BE",x"19C1",x"19C4",x"19C7",x"19CA",x"19CD",x"19D0",x"19D3",x"19D6",x"19D9",x"19DC",x"19DF",x"19E3",x"19E6",x"19E9",x"19EC",
x"19EF",x"19F2",x"19F5",x"19F8",x"19FB",x"19FE",x"1A01",x"1A04",x"1A07",x"1A0B",x"1A0E",x"1A11",x"1A14",x"1A17",x"1A1A",x"1A1D",
x"1A20",x"1A23",x"1A26",x"1A29",x"1A2C",x"1A2F",x"1A32",x"1A36",x"1A39",x"1A3C",x"1A3F",x"1A42",x"1A45",x"1A48",x"1A4B",x"1A4E",
x"1A51",x"1A54",x"1A57",x"1A5A",x"1A5E",x"1A61",x"1A64",x"1A67",x"1A6A",x"1A6D",x"1A70",x"1A73",x"1A76",x"1A79",x"1A7C",x"1A7F",
x"1A82",x"1A85",x"1A89",x"1A8C",x"1A8F",x"1A92",x"1A95",x"1A98",x"1A9B",x"1A9E",x"1AA1",x"1AA4",x"1AA7",x"1AAA",x"1AAD",x"1AB1",
x"1AB4",x"1AB7",x"1ABA",x"1ABD",x"1AC0",x"1AC3",x"1AC6",x"1AC9",x"1ACC",x"1ACF",x"1AD2",x"1AD5",x"1AD8",x"1ADC",x"1ADF",x"1AE2",
x"1AE5",x"1AE8",x"1AEB",x"1AEE",x"1AF1",x"1AF4",x"1AF7",x"1AFA",x"1AFD",x"1B00",x"1B03",x"1B07",x"1B0A",x"1B0D",x"1B10",x"1B13",
x"1B16",x"1B19",x"1B1C",x"1B1F",x"1B22",x"1B25",x"1B28",x"1B2B",x"1B2E",x"1B31",x"1B35",x"1B38",x"1B3B",x"1B3E",x"1B41",x"1B44",
x"1B47",x"1B4A",x"1B4D",x"1B50",x"1B53",x"1B56",x"1B59",x"1B5C",x"1B60",x"1B63",x"1B66",x"1B69",x"1B6C",x"1B6F",x"1B72",x"1B75",
x"1B78",x"1B7B",x"1B7E",x"1B81",x"1B84",x"1B87",x"1B8A",x"1B8E",x"1B91",x"1B94",x"1B97",x"1B9A",x"1B9D",x"1BA0",x"1BA3",x"1BA6",
x"1BA9",x"1BAC",x"1BAF",x"1BB2",x"1BB5",x"1BB9",x"1BBC",x"1BBF",x"1BC2",x"1BC5",x"1BC8",x"1BCB",x"1BCE",x"1BD1",x"1BD4",x"1BD7",
x"1BDA",x"1BDD",x"1BE0",x"1BE3",x"1BE7",x"1BEA",x"1BED",x"1BF0",x"1BF3",x"1BF6",x"1BF9",x"1BFC",x"1BFF",x"1C02",x"1C05",x"1C08",
x"1C0B",x"1C0E",x"1C11",x"1C14",x"1C18",x"1C1B",x"1C1E",x"1C21",x"1C24",x"1C27",x"1C2A",x"1C2D",x"1C30",x"1C33",x"1C36",x"1C39",
x"1C3C",x"1C3F",x"1C42",x"1C46",x"1C49",x"1C4C",x"1C4F",x"1C52",x"1C55",x"1C58",x"1C5B",x"1C5E",x"1C61",x"1C64",x"1C67",x"1C6A",
x"1C6D",x"1C70",x"1C73",x"1C77",x"1C7A",x"1C7D",x"1C80",x"1C83",x"1C86",x"1C89",x"1C8C",x"1C8F",x"1C92",x"1C95",x"1C98",x"1C9B",
x"1C9E",x"1CA1",x"1CA4",x"1CA8",x"1CAB",x"1CAE",x"1CB1",x"1CB4",x"1CB7",x"1CBA",x"1CBD",x"1CC0",x"1CC3",x"1CC6",x"1CC9",x"1CCC",
x"1CCF",x"1CD2",x"1CD5",x"1CD9",x"1CDC",x"1CDF",x"1CE2",x"1CE5",x"1CE8",x"1CEB",x"1CEE",x"1CF1",x"1CF4",x"1CF7",x"1CFA",x"1CFD",
x"1D00",x"1D03",x"1D06",x"1D09",x"1D0D",x"1D10",x"1D13",x"1D16",x"1D19",x"1D1C",x"1D1F",x"1D22",x"1D25",x"1D28",x"1D2B",x"1D2E",
x"1D31",x"1D34",x"1D37",x"1D3A",x"1D3D",x"1D41",x"1D44",x"1D47",x"1D4A",x"1D4D",x"1D50",x"1D53",x"1D56",x"1D59",x"1D5C",x"1D5F",
x"1D62",x"1D65",x"1D68",x"1D6B",x"1D6E",x"1D71",x"1D75",x"1D78",x"1D7B",x"1D7E",x"1D81",x"1D84",x"1D87",x"1D8A",x"1D8D",x"1D90",
x"1D93",x"1D96",x"1D99",x"1D9C",x"1D9F",x"1DA2",x"1DA5",x"1DA8",x"1DAC",x"1DAF",x"1DB2",x"1DB5",x"1DB8",x"1DBB",x"1DBE",x"1DC1",
x"1DC4",x"1DC7",x"1DCA",x"1DCD",x"1DD0",x"1DD3",x"1DD6",x"1DD9",x"1DDC",x"1DDF",x"1DE3",x"1DE6",x"1DE9",x"1DEC",x"1DEF",x"1DF2",
x"1DF5",x"1DF8",x"1DFB",x"1DFE",x"1E01",x"1E04",x"1E07",x"1E0A",x"1E0D",x"1E10",x"1E13",x"1E16",x"1E19",x"1E1D",x"1E20",x"1E23",
x"1E26",x"1E29",x"1E2C",x"1E2F",x"1E32",x"1E35",x"1E38",x"1E3B",x"1E3E",x"1E41",x"1E44",x"1E47",x"1E4A",x"1E4D",x"1E50",x"1E54",
x"1E57",x"1E5A",x"1E5D",x"1E60",x"1E63",x"1E66",x"1E69",x"1E6C",x"1E6F",x"1E72",x"1E75",x"1E78",x"1E7B",x"1E7E",x"1E81",x"1E84",
x"1E87",x"1E8A",x"1E8D",x"1E91",x"1E94",x"1E97",x"1E9A",x"1E9D",x"1EA0",x"1EA3",x"1EA6",x"1EA9",x"1EAC",x"1EAF",x"1EB2",x"1EB5",
x"1EB8",x"1EBB",x"1EBE",x"1EC1",x"1EC4",x"1EC7",x"1ECA",x"1ECE",x"1ED1",x"1ED4",x"1ED7",x"1EDA",x"1EDD",x"1EE0",x"1EE3",x"1EE6",
x"1EE9",x"1EEC",x"1EEF",x"1EF2",x"1EF5",x"1EF8",x"1EFB",x"1EFE",x"1F01",x"1F04",x"1F07",x"1F0A",x"1F0E",x"1F11",x"1F14",x"1F17",
x"1F1A",x"1F1D",x"1F20",x"1F23",x"1F26",x"1F29",x"1F2C",x"1F2F",x"1F32",x"1F35",x"1F38",x"1F3B",x"1F3E",x"1F41",x"1F44",x"1F47",
x"1F4A",x"1F4E",x"1F51",x"1F54",x"1F57",x"1F5A",x"1F5D",x"1F60",x"1F63",x"1F66",x"1F69",x"1F6C",x"1F6F",x"1F72",x"1F75",x"1F78",
x"1F7B",x"1F7E",x"1F81",x"1F84",x"1F87",x"1F8A",x"1F8D",x"1F91",x"1F94",x"1F97",x"1F9A",x"1F9D",x"1FA0",x"1FA3",x"1FA6",x"1FA9",
x"1FAC",x"1FAF",x"1FB2",x"1FB5",x"1FB8",x"1FBB",x"1FBE",x"1FC1",x"1FC4",x"1FC7",x"1FCA",x"1FCD",x"1FD0",x"1FD3",x"1FD7",x"1FDA",
x"1FDD",x"1FE0",x"1FE3",x"1FE6",x"1FE9",x"1FEC",x"1FEF",x"1FF2",x"1FF5",x"1FF8",x"1FFB",x"1FFE",x"2001",x"2004",x"2007",x"200A",
x"200D",x"2010",x"2013",x"2016",x"2019",x"201C",x"2020",x"2023",x"2026",x"2029",x"202C",x"202F",x"2032",x"2035",x"2038",x"203B",
x"203E",x"2041",x"2044",x"2047",x"204A",x"204D",x"2050",x"2053",x"2056",x"2059",x"205C",x"205F",x"2062",x"2065",x"2068",x"206C",
x"206F",x"2072",x"2075",x"2078",x"207B",x"207E",x"2081",x"2084",x"2087",x"208A",x"208D",x"2090",x"2093",x"2096",x"2099",x"209C",
x"209F",x"20A2",x"20A5",x"20A8",x"20AB",x"20AE",x"20B1",x"20B4",x"20B7",x"20BB",x"20BE",x"20C1",x"20C4",x"20C7",x"20CA",x"20CD",
x"20D0",x"20D3",x"20D6",x"20D9",x"20DC",x"20DF",x"20E2",x"20E5",x"20E8",x"20EB",x"20EE",x"20F1",x"20F4",x"20F7",x"20FA",x"20FD",
x"2100",x"2103",x"2106",x"2109",x"210C",x"2110",x"2113",x"2116",x"2119",x"211C",x"211F",x"2122",x"2125",x"2128",x"212B",x"212E",
x"2131",x"2134",x"2137",x"213A",x"213D",x"2140",x"2143",x"2146",x"2149",x"214C",x"214F",x"2152",x"2155",x"2158",x"215B",x"215E",
x"2161",x"2164",x"2168",x"216B",x"216E",x"2171",x"2174",x"2177",x"217A",x"217D",x"2180",x"2183",x"2186",x"2189",x"218C",x"218F",
x"2192",x"2195",x"2198",x"219B",x"219E",x"21A1",x"21A4",x"21A7",x"21AA",x"21AD",x"21B0",x"21B3",x"21B6",x"21B9",x"21BC",x"21BF",
x"21C2",x"21C5",x"21C9",x"21CC",x"21CF",x"21D2",x"21D5",x"21D8",x"21DB",x"21DE",x"21E1",x"21E4",x"21E7",x"21EA",x"21ED",x"21F0",
x"21F3",x"21F6",x"21F9",x"21FC",x"21FF",x"2202",x"2205",x"2208",x"220B",x"220E",x"2211",x"2214",x"2217",x"221A",x"221D",x"2220",
x"2223",x"2226",x"2229",x"222C",x"222F",x"2233",x"2236",x"2239",x"223C",x"223F",x"2242",x"2245",x"2248",x"224B",x"224E",x"2251",
x"2254",x"2257",x"225A",x"225D",x"2260",x"2263",x"2266",x"2269",x"226C",x"226F",x"2272",x"2275",x"2278",x"227B",x"227E",x"2281",
x"2284",x"2287",x"228A",x"228D",x"2290",x"2293",x"2296",x"2299",x"229C",x"229F",x"22A2",x"22A5",x"22A9",x"22AC",x"22AF",x"22B2",
x"22B5",x"22B8",x"22BB",x"22BE",x"22C1",x"22C4",x"22C7",x"22CA",x"22CD",x"22D0",x"22D3",x"22D6",x"22D9",x"22DC",x"22DF",x"22E2",
x"22E5",x"22E8",x"22EB",x"22EE",x"22F1",x"22F4",x"22F7",x"22FA",x"22FD",x"2300",x"2303",x"2306",x"2309",x"230C",x"230F",x"2312",
x"2315",x"2318",x"231B",x"231E",x"2321",x"2324",x"2327",x"232A",x"232E",x"2331",x"2334",x"2337",x"233A",x"233D",x"2340",x"2343",
x"2346",x"2349",x"234C",x"234F",x"2352",x"2355",x"2358",x"235B",x"235E",x"2361",x"2364",x"2367",x"236A",x"236D",x"2370",x"2373",
x"2376",x"2379",x"237C",x"237F",x"2382",x"2385",x"2388",x"238B",x"238E",x"2391",x"2394",x"2397",x"239A",x"239D",x"23A0",x"23A3",
x"23A6",x"23A9",x"23AC",x"23AF",x"23B2",x"23B5",x"23B8",x"23BB",x"23BE",x"23C1",x"23C4",x"23C7",x"23CA",x"23CD",x"23D0",x"23D4",
x"23D7",x"23DA",x"23DD",x"23E0",x"23E3",x"23E6",x"23E9",x"23EC",x"23EF",x"23F2",x"23F5",x"23F8",x"23FB",x"23FE",x"2401",x"2404",
x"2407",x"240A",x"240D",x"2410",x"2413",x"2416",x"2419",x"241C",x"241F",x"2422",x"2425",x"2428",x"242B",x"242E",x"2431",x"2434",
x"2437",x"243A",x"243D",x"2440",x"2443",x"2446",x"2449",x"244C",x"244F",x"2452",x"2455",x"2458",x"245B",x"245E",x"2461",x"2464",
x"2467",x"246A",x"246D",x"2470",x"2473",x"2476",x"2479",x"247C",x"247F",x"2482",x"2485",x"2488",x"248B",x"248E",x"2491",x"2494",
x"2497",x"249A",x"249D",x"24A0",x"24A3",x"24A6",x"24A9",x"24AC",x"24AF",x"24B2",x"24B5",x"24B8",x"24BB",x"24BE",x"24C1",x"24C5",
x"24C8",x"24CB",x"24CE",x"24D1",x"24D4",x"24D7",x"24DA",x"24DD",x"24E0",x"24E3",x"24E6",x"24E9",x"24EC",x"24EF",x"24F2",x"24F5",
x"24F8",x"24FB",x"24FE",x"2501",x"2504",x"2507",x"250A",x"250D",x"2510",x"2513",x"2516",x"2519",x"251C",x"251F",x"2522",x"2525",
x"2528",x"252B",x"252E",x"2531",x"2534",x"2537",x"253A",x"253D",x"2540",x"2543",x"2546",x"2549",x"254C",x"254F",x"2552",x"2555",
x"2558",x"255B",x"255E",x"2561",x"2564",x"2567",x"256A",x"256D",x"2570",x"2573",x"2576",x"2579",x"257C",x"257F",x"2582",x"2585",
x"2588",x"258B",x"258E",x"2591",x"2594",x"2597",x"259A",x"259D",x"25A0",x"25A3",x"25A6",x"25A9",x"25AC",x"25AF",x"25B2",x"25B5",
x"25B8",x"25BB",x"25BE",x"25C1",x"25C4",x"25C7",x"25CA",x"25CD",x"25D0",x"25D3",x"25D6",x"25D9",x"25DC",x"25DF",x"25E2",x"25E5",
x"25E8",x"25EB",x"25EE",x"25F1",x"25F4",x"25F7",x"25FA",x"25FD",x"2600",x"2603",x"2606",x"2609",x"260C",x"260F",x"2612",x"2615",
x"2618",x"261B",x"261E",x"2621",x"2624",x"2627",x"262A",x"262D",x"2630",x"2633",x"2636",x"2639",x"263C",x"263F",x"2642",x"2645",
x"2648",x"264B",x"264E",x"2651",x"2654",x"2657",x"265A",x"265D",x"2660",x"2663",x"2666",x"2669",x"266C",x"266F",x"2672",x"2675",
x"2678",x"267B",x"267E",x"2681",x"2684",x"2687",x"268A",x"268D",x"2690",x"2693",x"2696",x"2699",x"269C",x"269F",x"26A2",x"26A5",
x"26A8",x"26AB",x"26AE",x"26B1",x"26B4",x"26B7",x"26BA",x"26BD",x"26C0",x"26C3",x"26C6",x"26C9",x"26CC",x"26CF",x"26D2",x"26D5",
x"26D8",x"26DB",x"26DE",x"26E1",x"26E4",x"26E7",x"26EA",x"26ED",x"26F0",x"26F3",x"26F6",x"26F9",x"26FC",x"26FF",x"2702",x"2705",
x"2708",x"270B",x"270E",x"2711",x"2714",x"2717",x"271A",x"271D",x"2720",x"2723",x"2726",x"2729",x"272C",x"272F",x"2731",x"2734",
x"2737",x"273A",x"273D",x"2740",x"2743",x"2746",x"2749",x"274C",x"274F",x"2752",x"2755",x"2758",x"275B",x"275E",x"2761",x"2764",
x"2767",x"276A",x"276D",x"2770",x"2773",x"2776",x"2779",x"277C",x"277F",x"2782",x"2785",x"2788",x"278B",x"278E",x"2791",x"2794",
x"2797",x"279A",x"279D",x"27A0",x"27A3",x"27A6",x"27A9",x"27AC",x"27AF",x"27B2",x"27B5",x"27B8",x"27BB",x"27BE",x"27C1",x"27C4",
x"27C7",x"27CA",x"27CD",x"27D0",x"27D3",x"27D6",x"27D9",x"27DC",x"27DF",x"27E2",x"27E5",x"27E8",x"27EB",x"27EE",x"27F1",x"27F4",
x"27F7",x"27FA",x"27FD",x"2800",x"2803",x"2806",x"2809",x"280C",x"280F",x"2812",x"2815",x"2817",x"281A",x"281D",x"2820",x"2823",
x"2826",x"2829",x"282C",x"282F",x"2832",x"2835",x"2838",x"283B",x"283E",x"2841",x"2844",x"2847",x"284A",x"284D",x"2850",x"2853",
x"2856",x"2859",x"285C",x"285F",x"2862",x"2865",x"2868",x"286B",x"286E",x"2871",x"2874",x"2877",x"287A",x"287D",x"2880",x"2883",
x"2886",x"2889",x"288C",x"288F",x"2892",x"2895",x"2898",x"289B",x"289E",x"28A1",x"28A4",x"28A7",x"28AA",x"28AD",x"28B0",x"28B3",
x"28B5",x"28B8",x"28BB",x"28BE",x"28C1",x"28C4",x"28C7",x"28CA",x"28CD",x"28D0",x"28D3",x"28D6",x"28D9",x"28DC",x"28DF",x"28E2",
x"28E5",x"28E8",x"28EB",x"28EE",x"28F1",x"28F4",x"28F7",x"28FA",x"28FD",x"2900",x"2903",x"2906",x"2909",x"290C",x"290F",x"2912",
x"2915",x"2918",x"291B",x"291E",x"2921",x"2924",x"2927",x"292A",x"292D",x"2930",x"2932",x"2935",x"2938",x"293B",x"293E",x"2941",
x"2944",x"2947",x"294A",x"294D",x"2950",x"2953",x"2956",x"2959",x"295C",x"295F",x"2962",x"2965",x"2968",x"296B",x"296E",x"2971",
x"2974",x"2977",x"297A",x"297D",x"2980",x"2983",x"2986",x"2989",x"298C",x"298F",x"2992",x"2995",x"2998",x"299B",x"299E",x"29A0",
x"29A3",x"29A6",x"29A9",x"29AC",x"29AF",x"29B2",x"29B5",x"29B8",x"29BB",x"29BE",x"29C1",x"29C4",x"29C7",x"29CA",x"29CD",x"29D0",
x"29D3",x"29D6",x"29D9",x"29DC",x"29DF",x"29E2",x"29E5",x"29E8",x"29EB",x"29EE",x"29F1",x"29F4",x"29F7",x"29FA",x"29FD",x"29FF",
x"2A02",x"2A05",x"2A08",x"2A0B",x"2A0E",x"2A11",x"2A14",x"2A17",x"2A1A",x"2A1D",x"2A20",x"2A23",x"2A26",x"2A29",x"2A2C",x"2A2F",
x"2A32",x"2A35",x"2A38",x"2A3B",x"2A3E",x"2A41",x"2A44",x"2A47",x"2A4A",x"2A4D",x"2A50",x"2A53",x"2A56",x"2A58",x"2A5B",x"2A5E",
x"2A61",x"2A64",x"2A67",x"2A6A",x"2A6D",x"2A70",x"2A73",x"2A76",x"2A79",x"2A7C",x"2A7F",x"2A82",x"2A85",x"2A88",x"2A8B",x"2A8E",
x"2A91",x"2A94",x"2A97",x"2A9A",x"2A9D",x"2AA0",x"2AA3",x"2AA6",x"2AA8",x"2AAB",x"2AAE",x"2AB1",x"2AB4",x"2AB7",x"2ABA",x"2ABD",
x"2AC0",x"2AC3",x"2AC6",x"2AC9",x"2ACC",x"2ACF",x"2AD2",x"2AD5",x"2AD8",x"2ADB",x"2ADE",x"2AE1",x"2AE4",x"2AE7",x"2AEA",x"2AED",
x"2AF0",x"2AF2",x"2AF5",x"2AF8",x"2AFB",x"2AFE",x"2B01",x"2B04",x"2B07",x"2B0A",x"2B0D",x"2B10",x"2B13",x"2B16",x"2B19",x"2B1C",
x"2B1F",x"2B22",x"2B25",x"2B28",x"2B2B",x"2B2E",x"2B31",x"2B34",x"2B37",x"2B39",x"2B3C",x"2B3F",x"2B42",x"2B45",x"2B48",x"2B4B",
x"2B4E",x"2B51",x"2B54",x"2B57",x"2B5A",x"2B5D",x"2B60",x"2B63",x"2B66",x"2B69",x"2B6C",x"2B6F",x"2B72",x"2B75",x"2B78",x"2B7B",
x"2B7D",x"2B80",x"2B83",x"2B86",x"2B89",x"2B8C",x"2B8F",x"2B92",x"2B95",x"2B98",x"2B9B",x"2B9E",x"2BA1",x"2BA4",x"2BA7",x"2BAA",
x"2BAD",x"2BB0",x"2BB3",x"2BB6",x"2BB9",x"2BBB",x"2BBE",x"2BC1",x"2BC4",x"2BC7",x"2BCA",x"2BCD",x"2BD0",x"2BD3",x"2BD6",x"2BD9",
x"2BDC",x"2BDF",x"2BE2",x"2BE5",x"2BE8",x"2BEB",x"2BEE",x"2BF1",x"2BF4",x"2BF7",x"2BF9",x"2BFC",x"2BFF",x"2C02",x"2C05",x"2C08",
x"2C0B",x"2C0E",x"2C11",x"2C14",x"2C17",x"2C1A",x"2C1D",x"2C20",x"2C23",x"2C26",x"2C29",x"2C2C",x"2C2F",x"2C32",x"2C34",x"2C37",
x"2C3A",x"2C3D",x"2C40",x"2C43",x"2C46",x"2C49",x"2C4C",x"2C4F",x"2C52",x"2C55",x"2C58",x"2C5B",x"2C5E",x"2C61",x"2C64",x"2C67",
x"2C6A",x"2C6C",x"2C6F",x"2C72",x"2C75",x"2C78",x"2C7B",x"2C7E",x"2C81",x"2C84",x"2C87",x"2C8A",x"2C8D",x"2C90",x"2C93",x"2C96",
x"2C99",x"2C9C",x"2C9F",x"2CA1",x"2CA4",x"2CA7",x"2CAA",x"2CAD",x"2CB0",x"2CB3",x"2CB6",x"2CB9",x"2CBC",x"2CBF",x"2CC2",x"2CC5",
x"2CC8",x"2CCB",x"2CCE",x"2CD1",x"2CD4",x"2CD6",x"2CD9",x"2CDC",x"2CDF",x"2CE2",x"2CE5",x"2CE8",x"2CEB",x"2CEE",x"2CF1",x"2CF4",
x"2CF7",x"2CFA",x"2CFD",x"2D00",x"2D03",x"2D06",x"2D08",x"2D0B",x"2D0E",x"2D11",x"2D14",x"2D17",x"2D1A",x"2D1D",x"2D20",x"2D23",
x"2D26",x"2D29",x"2D2C",x"2D2F",x"2D32",x"2D35",x"2D37",x"2D3A",x"2D3D",x"2D40",x"2D43",x"2D46",x"2D49",x"2D4C",x"2D4F",x"2D52",
x"2D55",x"2D58",x"2D5B",x"2D5E",x"2D61",x"2D64",x"2D67",x"2D69",x"2D6C",x"2D6F",x"2D72",x"2D75",x"2D78",x"2D7B",x"2D7E",x"2D81",
x"2D84",x"2D87",x"2D8A",x"2D8D",x"2D90",x"2D93",x"2D95",x"2D98",x"2D9B",x"2D9E",x"2DA1",x"2DA4",x"2DA7",x"2DAA",x"2DAD",x"2DB0",
x"2DB3",x"2DB6",x"2DB9",x"2DBC",x"2DBF",x"2DC2",x"2DC4",x"2DC7",x"2DCA",x"2DCD",x"2DD0",x"2DD3",x"2DD6",x"2DD9",x"2DDC",x"2DDF",
x"2DE2",x"2DE5",x"2DE8",x"2DEB",x"2DEE",x"2DF0",x"2DF3",x"2DF6",x"2DF9",x"2DFC",x"2DFF",x"2E02",x"2E05",x"2E08",x"2E0B",x"2E0E",
x"2E11",x"2E14",x"2E17",x"2E19",x"2E1C",x"2E1F",x"2E22",x"2E25",x"2E28",x"2E2B",x"2E2E",x"2E31",x"2E34",x"2E37",x"2E3A",x"2E3D",
x"2E40",x"2E42",x"2E45",x"2E48",x"2E4B",x"2E4E",x"2E51",x"2E54",x"2E57",x"2E5A",x"2E5D",x"2E60",x"2E63",x"2E66",x"2E69",x"2E6B",
x"2E6E",x"2E71",x"2E74",x"2E77",x"2E7A",x"2E7D",x"2E80",x"2E83",x"2E86",x"2E89",x"2E8C",x"2E8F",x"2E92",x"2E94",x"2E97",x"2E9A",
x"2E9D",x"2EA0",x"2EA3",x"2EA6",x"2EA9",x"2EAC",x"2EAF",x"2EB2",x"2EB5",x"2EB8",x"2EBA",x"2EBD",x"2EC0",x"2EC3",x"2EC6",x"2EC9",
x"2ECC",x"2ECF",x"2ED2",x"2ED5",x"2ED8",x"2EDB",x"2EDE",x"2EE1",x"2EE3",x"2EE6",x"2EE9",x"2EEC",x"2EEF",x"2EF2",x"2EF5",x"2EF8",
x"2EFB",x"2EFE",x"2F01",x"2F04",x"2F06",x"2F09",x"2F0C",x"2F0F",x"2F12",x"2F15",x"2F18",x"2F1B",x"2F1E",x"2F21",x"2F24",x"2F27",
x"2F2A",x"2F2C",x"2F2F",x"2F32",x"2F35",x"2F38",x"2F3B",x"2F3E",x"2F41",x"2F44",x"2F47",x"2F4A",x"2F4D",x"2F50",x"2F52",x"2F55",
x"2F58",x"2F5B",x"2F5E",x"2F61",x"2F64",x"2F67",x"2F6A",x"2F6D",x"2F70",x"2F73",x"2F75",x"2F78",x"2F7B",x"2F7E",x"2F81",x"2F84",
x"2F87",x"2F8A",x"2F8D",x"2F90",x"2F93",x"2F96",x"2F98",x"2F9B",x"2F9E",x"2FA1",x"2FA4",x"2FA7",x"2FAA",x"2FAD",x"2FB0",x"2FB3",
x"2FB6",x"2FB9",x"2FBB",x"2FBE",x"2FC1",x"2FC4",x"2FC7",x"2FCA",x"2FCD",x"2FD0",x"2FD3",x"2FD6",x"2FD9",x"2FDB",x"2FDE",x"2FE1",
x"2FE4",x"2FE7",x"2FEA",x"2FED",x"2FF0",x"2FF3",x"2FF6",x"2FF9",x"2FFC",x"2FFE",x"3001",x"3004",x"3007",x"300A",x"300D",x"3010",
x"3013",x"3016",x"3019",x"301C",x"301E",x"3021",x"3024",x"3027",x"302A",x"302D",x"3030",x"3033",x"3036",x"3039",x"303C",x"303E",
x"3041",x"3044",x"3047",x"304A",x"304D",x"3050",x"3053",x"3056",x"3059",x"305C",x"305E",x"3061",x"3064",x"3067",x"306A",x"306D",
x"3070",x"3073",x"3076",x"3079",x"307C",x"307E",x"3081",x"3084",x"3087",x"308A",x"308D",x"3090",x"3093",x"3096",x"3099",x"309C",
x"309E",x"30A1",x"30A4",x"30A7",x"30AA",x"30AD",x"30B0",x"30B3",x"30B6",x"30B9",x"30BC",x"30BE",x"30C1",x"30C4",x"30C7",x"30CA",
x"30CD",x"30D0",x"30D3",x"30D6",x"30D9",x"30DB",x"30DE",x"30E1",x"30E4",x"30E7",x"30EA",x"30ED",x"30F0",x"30F3",x"30F6",x"30F8",
x"30FB",x"30FE",x"3101",x"3104",x"3107",x"310A",x"310D",x"3110",x"3113",x"3116",x"3118",x"311B",x"311E",x"3121",x"3124",x"3127",
x"312A",x"312D",x"3130",x"3133",x"3135",x"3138",x"313B",x"313E",x"3141",x"3144",x"3147",x"314A",x"314D",x"3150",x"3152",x"3155",
x"3158",x"315B",x"315E",x"3161",x"3164",x"3167",x"316A",x"316C",x"316F",x"3172",x"3175",x"3178",x"317B",x"317E",x"3181",x"3184",
x"3187",x"3189",x"318C",x"318F",x"3192",x"3195",x"3198",x"319B",x"319E",x"31A1",x"31A4",x"31A6",x"31A9",x"31AC",x"31AF",x"31B2",
x"31B5",x"31B8",x"31BB",x"31BE",x"31C0",x"31C3",x"31C6",x"31C9",x"31CC",x"31CF",x"31D2",x"31D5",x"31D8",x"31DB",x"31DD",x"31E0",
x"31E3",x"31E6",x"31E9",x"31EC",x"31EF",x"31F2",x"31F5",x"31F7",x"31FA",x"31FD",x"3200",x"3203",x"3206",x"3209",x"320C",x"320F",
x"3211",x"3214",x"3217",x"321A",x"321D",x"3220",x"3223",x"3226",x"3229",x"322B",x"322E",x"3231",x"3234",x"3237",x"323A",x"323D",
x"3240",x"3243",x"3246",x"3248",x"324B",x"324E",x"3251",x"3254",x"3257",x"325A",x"325D",x"325F",x"3262",x"3265",x"3268",x"326B",
x"326E",x"3271",x"3274",x"3277",x"3279",x"327C",x"327F",x"3282",x"3285",x"3288",x"328B",x"328E",x"3291",x"3293",x"3296",x"3299",
x"329C",x"329F",x"32A2",x"32A5",x"32A8",x"32AB",x"32AD",x"32B0",x"32B3",x"32B6",x"32B9",x"32BC",x"32BF",x"32C2",x"32C5",x"32C7",
x"32CA",x"32CD",x"32D0",x"32D3",x"32D6",x"32D9",x"32DC",x"32DE",x"32E1",x"32E4",x"32E7",x"32EA",x"32ED",x"32F0",x"32F3",x"32F6",
x"32F8",x"32FB",x"32FE",x"3301",x"3304",x"3307",x"330A",x"330D",x"330F",x"3312",x"3315",x"3318",x"331B",x"331E",x"3321",x"3324",
x"3326",x"3329",x"332C",x"332F",x"3332",x"3335",x"3338",x"333B",x"333E",x"3340",x"3343",x"3346",x"3349",x"334C",x"334F",x"3352",
x"3355",x"3357",x"335A",x"335D",x"3360",x"3363",x"3366",x"3369",x"336C",x"336E",x"3371",x"3374",x"3377",x"337A",x"337D",x"3380",
x"3383",x"3385",x"3388",x"338B",x"338E",x"3391",x"3394",x"3397",x"339A",x"339C",x"339F",x"33A2",x"33A5",x"33A8",x"33AB",x"33AE",
x"33B1",x"33B3",x"33B6",x"33B9",x"33BC",x"33BF",x"33C2",x"33C5",x"33C8",x"33CA",x"33CD",x"33D0",x"33D3",x"33D6",x"33D9",x"33DC",
x"33DF",x"33E1",x"33E4",x"33E7",x"33EA",x"33ED",x"33F0",x"33F3",x"33F6",x"33F8",x"33FB",x"33FE",x"3401",x"3404",x"3407",x"340A",
x"340C",x"340F",x"3412",x"3415",x"3418",x"341B",x"341E",x"3421",x"3423",x"3426",x"3429",x"342C",x"342F",x"3432",x"3435",x"3438",
x"343A",x"343D",x"3440",x"3443",x"3446",x"3449",x"344C",x"344E",x"3451",x"3454",x"3457",x"345A",x"345D",x"3460",x"3463",x"3465",
x"3468",x"346B",x"346E",x"3471",x"3474",x"3477",x"3479",x"347C",x"347F",x"3482",x"3485",x"3488",x"348B",x"348E",x"3490",x"3493",
x"3496",x"3499",x"349C",x"349F",x"34A2",x"34A4",x"34A7",x"34AA",x"34AD",x"34B0",x"34B3",x"34B6",x"34B8",x"34BB",x"34BE",x"34C1",
x"34C4",x"34C7",x"34CA",x"34CC",x"34CF",x"34D2",x"34D5",x"34D8",x"34DB",x"34DE",x"34E1",x"34E3",x"34E6",x"34E9",x"34EC",x"34EF",
x"34F2",x"34F5",x"34F7",x"34FA",x"34FD",x"3500",x"3503",x"3506",x"3509",x"350B",x"350E",x"3511",x"3514",x"3517",x"351A",x"351D",
x"351F",x"3522",x"3525",x"3528",x"352B",x"352E",x"3531",x"3533",x"3536",x"3539",x"353C",x"353F",x"3542",x"3545",x"3547",x"354A",
x"354D",x"3550",x"3553",x"3556",x"3559",x"355B",x"355E",x"3561",x"3564",x"3567",x"356A",x"356D",x"356F",x"3572",x"3575",x"3578",
x"357B",x"357E",x"3581",x"3583",x"3586",x"3589",x"358C",x"358F",x"3592",x"3595",x"3597",x"359A",x"359D",x"35A0",x"35A3",x"35A6",
x"35A8",x"35AB",x"35AE",x"35B1",x"35B4",x"35B7",x"35BA",x"35BC",x"35BF",x"35C2",x"35C5",x"35C8",x"35CB",x"35CE",x"35D0",x"35D3",
x"35D6",x"35D9",x"35DC",x"35DF",x"35E1",x"35E4",x"35E7",x"35EA",x"35ED",x"35F0",x"35F3",x"35F5",x"35F8",x"35FB",x"35FE",x"3601",
x"3604",x"3607",x"3609",x"360C",x"360F",x"3612",x"3615",x"3618",x"361A",x"361D",x"3620",x"3623",x"3626",x"3629",x"362C",x"362E",
x"3631",x"3634",x"3637",x"363A",x"363D",x"363F",x"3642",x"3645",x"3648",x"364B",x"364E",x"3651",x"3653",x"3656",x"3659",x"365C",
x"365F",x"3662",x"3664",x"3667",x"366A",x"366D",x"3670",x"3673",x"3676",x"3678",x"367B",x"367E",x"3681",x"3684",x"3687",x"3689",
x"368C",x"368F",x"3692",x"3695",x"3698",x"369A",x"369D",x"36A0",x"36A3",x"36A6",x"36A9",x"36AB",x"36AE",x"36B1",x"36B4",x"36B7",
x"36BA",x"36BD",x"36BF",x"36C2",x"36C5",x"36C8",x"36CB",x"36CE",x"36D0",x"36D3",x"36D6",x"36D9",x"36DC",x"36DF",x"36E1",x"36E4",
x"36E7",x"36EA",x"36ED",x"36F0",x"36F2",x"36F5",x"36F8",x"36FB",x"36FE",x"3701",x"3703",x"3706",x"3709",x"370C",x"370F",x"3712",
x"3715",x"3717",x"371A",x"371D",x"3720",x"3723",x"3726",x"3728",x"372B",x"372E",x"3731",x"3734",x"3737",x"3739",x"373C",x"373F",
x"3742",x"3745",x"3748",x"374A",x"374D",x"3750",x"3753",x"3756",x"3759",x"375B",x"375E",x"3761",x"3764",x"3767",x"376A",x"376C",
x"376F",x"3772",x"3775",x"3778",x"377B",x"377D",x"3780",x"3783",x"3786",x"3789",x"378B",x"378E",x"3791",x"3794",x"3797",x"379A",
x"379C",x"379F",x"37A2",x"37A5",x"37A8",x"37AB",x"37AD",x"37B0",x"37B3",x"37B6",x"37B9",x"37BC",x"37BE",x"37C1",x"37C4",x"37C7",
x"37CA",x"37CD",x"37CF",x"37D2",x"37D5",x"37D8",x"37DB",x"37DE",x"37E0",x"37E3",x"37E6",x"37E9",x"37EC",x"37EE",x"37F1",x"37F4",
x"37F7",x"37FA",x"37FD",x"37FF",x"3802",x"3805",x"3808",x"380B",x"380E",x"3810",x"3813",x"3816",x"3819",x"381C",x"381E",x"3821",
x"3824",x"3827",x"382A",x"382D",x"382F",x"3832",x"3835",x"3838",x"383B",x"383E",x"3840",x"3843",x"3846",x"3849",x"384C",x"384E",
x"3851",x"3854",x"3857",x"385A",x"385D",x"385F",x"3862",x"3865",x"3868",x"386B",x"386D",x"3870",x"3873",x"3876",x"3879",x"387C",
x"387E",x"3881",x"3884",x"3887",x"388A",x"388D",x"388F",x"3892",x"3895",x"3898",x"389B",x"389D",x"38A0",x"38A3",x"38A6",x"38A9",
x"38AB",x"38AE",x"38B1",x"38B4",x"38B7",x"38BA",x"38BC",x"38BF",x"38C2",x"38C5",x"38C8",x"38CA",x"38CD",x"38D0",x"38D3",x"38D6",
x"38D9",x"38DB",x"38DE",x"38E1",x"38E4",x"38E7",x"38E9",x"38EC",x"38EF",x"38F2",x"38F5",x"38F8",x"38FA",x"38FD",x"3900",x"3903",
x"3906",x"3908",x"390B",x"390E",x"3911",x"3914",x"3916",x"3919",x"391C",x"391F",x"3922",x"3924",x"3927",x"392A",x"392D",x"3930",
x"3933",x"3935",x"3938",x"393B",x"393E",x"3941",x"3943",x"3946",x"3949",x"394C",x"394F",x"3951",x"3954",x"3957",x"395A",x"395D",
x"3960",x"3962",x"3965",x"3968",x"396B",x"396E",x"3970",x"3973",x"3976",x"3979",x"397C",x"397E",x"3981",x"3984",x"3987",x"398A",
x"398C",x"398F",x"3992",x"3995",x"3998",x"399A",x"399D",x"39A0",x"39A3",x"39A6",x"39A8",x"39AB",x"39AE",x"39B1",x"39B4",x"39B6",
x"39B9",x"39BC",x"39BF",x"39C2",x"39C5",x"39C7",x"39CA",x"39CD",x"39D0",x"39D3",x"39D5",x"39D8",x"39DB",x"39DE",x"39E1",x"39E3",
x"39E6",x"39E9",x"39EC",x"39EF",x"39F1",x"39F4",x"39F7",x"39FA",x"39FD",x"39FF",x"3A02",x"3A05",x"3A08",x"3A0B",x"3A0D",x"3A10",
x"3A13",x"3A16",x"3A19",x"3A1B",x"3A1E",x"3A21",x"3A24",x"3A27",x"3A29",x"3A2C",x"3A2F",x"3A32",x"3A35",x"3A37",x"3A3A",x"3A3D",
x"3A40",x"3A43",x"3A45",x"3A48",x"3A4B",x"3A4E",x"3A51",x"3A53",x"3A56",x"3A59",x"3A5C",x"3A5E",x"3A61",x"3A64",x"3A67",x"3A6A",
x"3A6C",x"3A6F",x"3A72",x"3A75",x"3A78",x"3A7A",x"3A7D",x"3A80",x"3A83",x"3A86",x"3A88",x"3A8B",x"3A8E",x"3A91",x"3A94",x"3A96",
x"3A99",x"3A9C",x"3A9F",x"3AA2",x"3AA4",x"3AA7",x"3AAA",x"3AAD",x"3AB0",x"3AB2",x"3AB5",x"3AB8",x"3ABB",x"3ABD",x"3AC0",x"3AC3",
x"3AC6",x"3AC9",x"3ACB",x"3ACE",x"3AD1",x"3AD4",x"3AD7",x"3AD9",x"3ADC",x"3ADF",x"3AE2",x"3AE5",x"3AE7",x"3AEA",x"3AED",x"3AF0",
x"3AF2",x"3AF5",x"3AF8",x"3AFB",x"3AFE",x"3B00",x"3B03",x"3B06",x"3B09",x"3B0C",x"3B0E",x"3B11",x"3B14",x"3B17",x"3B19",x"3B1C",
x"3B1F",x"3B22",x"3B25",x"3B27",x"3B2A",x"3B2D",x"3B30",x"3B33",x"3B35",x"3B38",x"3B3B",x"3B3E",x"3B40",x"3B43",x"3B46",x"3B49",
x"3B4C",x"3B4E",x"3B51",x"3B54",x"3B57",x"3B5A",x"3B5C",x"3B5F",x"3B62",x"3B65",x"3B67",x"3B6A",x"3B6D",x"3B70",x"3B73",x"3B75",
x"3B78",x"3B7B",x"3B7E",x"3B81",x"3B83",x"3B86",x"3B89",x"3B8C",x"3B8E",x"3B91",x"3B94",x"3B97",x"3B9A",x"3B9C",x"3B9F",x"3BA2",
x"3BA5",x"3BA7",x"3BAA",x"3BAD",x"3BB0",x"3BB3",x"3BB5",x"3BB8",x"3BBB",x"3BBE",x"3BC0",x"3BC3",x"3BC6",x"3BC9",x"3BCC",x"3BCE",
x"3BD1",x"3BD4",x"3BD7",x"3BD9",x"3BDC",x"3BDF",x"3BE2",x"3BE5",x"3BE7",x"3BEA",x"3BED",x"3BF0",x"3BF2",x"3BF5",x"3BF8",x"3BFB",
x"3BFE",x"3C00",x"3C03",x"3C06",x"3C09",x"3C0B",x"3C0E",x"3C11",x"3C14",x"3C16",x"3C19",x"3C1C",x"3C1F",x"3C22",x"3C24",x"3C27",
x"3C2A",x"3C2D",x"3C2F",x"3C32",x"3C35",x"3C38",x"3C3B",x"3C3D",x"3C40",x"3C43",x"3C46",x"3C48",x"3C4B",x"3C4E",x"3C51",x"3C53",
x"3C56",x"3C59",x"3C5C",x"3C5F",x"3C61",x"3C64",x"3C67",x"3C6A",x"3C6C",x"3C6F",x"3C72",x"3C75",x"3C77",x"3C7A",x"3C7D",x"3C80",
x"3C83",x"3C85",x"3C88",x"3C8B",x"3C8E",x"3C90",x"3C93",x"3C96",x"3C99",x"3C9B",x"3C9E",x"3CA1",x"3CA4",x"3CA7",x"3CA9",x"3CAC",
x"3CAF",x"3CB2",x"3CB4",x"3CB7",x"3CBA",x"3CBD",x"3CBF",x"3CC2",x"3CC5",x"3CC8",x"3CCA",x"3CCD",x"3CD0",x"3CD3",x"3CD6",x"3CD8",
x"3CDB",x"3CDE",x"3CE1",x"3CE3",x"3CE6",x"3CE9",x"3CEC",x"3CEE",x"3CF1",x"3CF4",x"3CF7",x"3CF9",x"3CFC",x"3CFF",x"3D02",x"3D05",
x"3D07",x"3D0A",x"3D0D",x"3D10",x"3D12",x"3D15",x"3D18",x"3D1B",x"3D1D",x"3D20",x"3D23",x"3D26",x"3D28",x"3D2B",x"3D2E",x"3D31",
x"3D33",x"3D36",x"3D39",x"3D3C",x"3D3E",x"3D41",x"3D44",x"3D47",x"3D4A",x"3D4C",x"3D4F",x"3D52",x"3D55",x"3D57",x"3D5A",x"3D5D",
x"3D60",x"3D62",x"3D65",x"3D68",x"3D6B",x"3D6D",x"3D70",x"3D73",x"3D76",x"3D78",x"3D7B",x"3D7E",x"3D81",x"3D83",x"3D86",x"3D89",
x"3D8C",x"3D8E",x"3D91",x"3D94",x"3D97",x"3D99",x"3D9C",x"3D9F",x"3DA2",x"3DA4",x"3DA7",x"3DAA",x"3DAD",x"3DAF",x"3DB2",x"3DB5",
x"3DB8",x"3DBA",x"3DBD",x"3DC0",x"3DC3",x"3DC5",x"3DC8",x"3DCB",x"3DCE",x"3DD0",x"3DD3",x"3DD6",x"3DD9",x"3DDB",x"3DDE",x"3DE1",
x"3DE4",x"3DE6",x"3DE9",x"3DEC",x"3DEF",x"3DF1",x"3DF4",x"3DF7",x"3DFA",x"3DFC",x"3DFF",x"3E02",x"3E05",x"3E07",x"3E0A",x"3E0D",
x"3E10",x"3E12",x"3E15",x"3E18",x"3E1B",x"3E1D",x"3E20",x"3E23",x"3E26",x"3E28",x"3E2B",x"3E2E",x"3E31",x"3E33",x"3E36",x"3E39",
x"3E3C",x"3E3E",x"3E41",x"3E44",x"3E47",x"3E49",x"3E4C",x"3E4F",x"3E52",x"3E54",x"3E57",x"3E5A",x"3E5D",x"3E5F",x"3E62",x"3E65",
x"3E68",x"3E6A",x"3E6D",x"3E70",x"3E73",x"3E75",x"3E78",x"3E7B",x"3E7D",x"3E80",x"3E83",x"3E86",x"3E88",x"3E8B",x"3E8E",x"3E91",
x"3E93",x"3E96",x"3E99",x"3E9C",x"3E9E",x"3EA1",x"3EA4",x"3EA7",x"3EA9",x"3EAC",x"3EAF",x"3EB2",x"3EB4",x"3EB7",x"3EBA",x"3EBD",
x"3EBF",x"3EC2",x"3EC5",x"3EC7",x"3ECA",x"3ECD",x"3ED0",x"3ED2",x"3ED5",x"3ED8",x"3EDB",x"3EDD",x"3EE0",x"3EE3",x"3EE6",x"3EE8",
x"3EEB",x"3EEE",x"3EF1",x"3EF3",x"3EF6",x"3EF9",x"3EFB",x"3EFE",x"3F01",x"3F04",x"3F06",x"3F09",x"3F0C",x"3F0F",x"3F11",x"3F14",
x"3F17",x"3F1A",x"3F1C",x"3F1F",x"3F22",x"3F24",x"3F27",x"3F2A",x"3F2D",x"3F2F",x"3F32",x"3F35",x"3F38",x"3F3A",x"3F3D",x"3F40",
x"3F43",x"3F45",x"3F48",x"3F4B",x"3F4D",x"3F50",x"3F53",x"3F56",x"3F58",x"3F5B",x"3F5E",x"3F61",x"3F63",x"3F66",x"3F69",x"3F6B",
x"3F6E",x"3F71",x"3F74",x"3F76",x"3F79",x"3F7C",x"3F7F",x"3F81",x"3F84",x"3F87",x"3F89",x"3F8C",x"3F8F",x"3F92",x"3F94",x"3F97",
x"3F9A",x"3F9D",x"3F9F",x"3FA2",x"3FA5",x"3FA7",x"3FAA",x"3FAD",x"3FB0",x"3FB2",x"3FB5",x"3FB8",x"3FBB",x"3FBD",x"3FC0",x"3FC3",
x"3FC5",x"3FC8",x"3FCB",x"3FCE",x"3FD0",x"3FD3",x"3FD6",x"3FD8",x"3FDB",x"3FDE",x"3FE1",x"3FE3",x"3FE6",x"3FE9",x"3FEC",x"3FEE",
x"3FF1",x"3FF4",x"3FF6",x"3FF9",x"3FFC",x"3FFF",x"4001",x"4004",x"4007",x"4009",x"400C",x"400F",x"4012",x"4014",x"4017",x"401A",
x"401D",x"401F",x"4022",x"4025",x"4027",x"402A",x"402D",x"4030",x"4032",x"4035",x"4038",x"403A",x"403D",x"4040",x"4043",x"4045",
x"4048",x"404B",x"404D",x"4050",x"4053",x"4056",x"4058",x"405B",x"405E",x"4060",x"4063",x"4066",x"4069",x"406B",x"406E",x"4071",
x"4073",x"4076",x"4079",x"407C",x"407E",x"4081",x"4084",x"4086",x"4089",x"408C",x"408F",x"4091",x"4094",x"4097",x"4099",x"409C",
x"409F",x"40A2",x"40A4",x"40A7",x"40AA",x"40AC",x"40AF",x"40B2",x"40B5",x"40B7",x"40BA",x"40BD",x"40BF",x"40C2",x"40C5",x"40C8",
x"40CA",x"40CD",x"40D0",x"40D2",x"40D5",x"40D8",x"40DA",x"40DD",x"40E0",x"40E3",x"40E5",x"40E8",x"40EB",x"40ED",x"40F0",x"40F3",
x"40F6",x"40F8",x"40FB",x"40FE",x"4100",x"4103",x"4106",x"4108",x"410B",x"410E",x"4111",x"4113",x"4116",x"4119",x"411B",x"411E",
x"4121",x"4124",x"4126",x"4129",x"412C",x"412E",x"4131",x"4134",x"4136",x"4139",x"413C",x"413F",x"4141",x"4144",x"4147",x"4149",
x"414C",x"414F",x"4151",x"4154",x"4157",x"415A",x"415C",x"415F",x"4162",x"4164",x"4167",x"416A",x"416D",x"416F",x"4172",x"4175",
x"4177",x"417A",x"417D",x"417F",x"4182",x"4185",x"4187",x"418A",x"418D",x"4190",x"4192",x"4195",x"4198",x"419A",x"419D",x"41A0",
x"41A2",x"41A5",x"41A8",x"41AB",x"41AD",x"41B0",x"41B3",x"41B5",x"41B8",x"41BB",x"41BD",x"41C0",x"41C3",x"41C6",x"41C8",x"41CB",
x"41CE",x"41D0",x"41D3",x"41D6",x"41D8",x"41DB",x"41DE",x"41E0",x"41E3",x"41E6",x"41E9",x"41EB",x"41EE",x"41F1",x"41F3",x"41F6",
x"41F9",x"41FB",x"41FE",x"4201",x"4203",x"4206",x"4209",x"420C",x"420E",x"4211",x"4214",x"4216",x"4219",x"421C",x"421E",x"4221",
x"4224",x"4226",x"4229",x"422C",x"422F",x"4231",x"4234",x"4237",x"4239",x"423C",x"423F",x"4241",x"4244",x"4247",x"4249",x"424C",
x"424F",x"4251",x"4254",x"4257",x"425A",x"425C",x"425F",x"4262",x"4264",x"4267",x"426A",x"426C",x"426F",x"4272",x"4274",x"4277",
x"427A",x"427C",x"427F",x"4282",x"4284",x"4287",x"428A",x"428D",x"428F",x"4292",x"4295",x"4297",x"429A",x"429D",x"429F",x"42A2",
x"42A5",x"42A7",x"42AA",x"42AD",x"42AF",x"42B2",x"42B5",x"42B7",x"42BA",x"42BD",x"42BF",x"42C2",x"42C5",x"42C8",x"42CA",x"42CD",
x"42D0",x"42D2",x"42D5",x"42D8",x"42DA",x"42DD",x"42E0",x"42E2",x"42E5",x"42E8",x"42EA",x"42ED",x"42F0",x"42F2",x"42F5",x"42F8",
x"42FA",x"42FD",x"4300",x"4302",x"4305",x"4308",x"430A",x"430D",x"4310",x"4313",x"4315",x"4318",x"431B",x"431D",x"4320",x"4323",
x"4325",x"4328",x"432B",x"432D",x"4330",x"4333",x"4335",x"4338",x"433B",x"433D",x"4340",x"4343",x"4345",x"4348",x"434B",x"434D",
x"4350",x"4353",x"4355",x"4358",x"435B",x"435D",x"4360",x"4363",x"4365",x"4368",x"436B",x"436D",x"4370",x"4373",x"4375",x"4378",
x"437B",x"437D",x"4380",x"4383",x"4385",x"4388",x"438B",x"438D",x"4390",x"4393",x"4395",x"4398",x"439B",x"439D",x"43A0",x"43A3",
x"43A5",x"43A8",x"43AB",x"43AD",x"43B0",x"43B3",x"43B5",x"43B8",x"43BB",x"43BD",x"43C0",x"43C3",x"43C5",x"43C8",x"43CB",x"43CD",
x"43D0",x"43D3",x"43D5",x"43D8",x"43DB",x"43DD",x"43E0",x"43E3",x"43E5",x"43E8",x"43EB",x"43ED",x"43F0",x"43F3",x"43F5",x"43F8",
x"43FB",x"43FD",x"4400",x"4403",x"4405",x"4408",x"440B",x"440D",x"4410",x"4413",x"4415",x"4418",x"441B",x"441D",x"4420",x"4423",
x"4425",x"4428",x"442B",x"442D",x"4430",x"4433",x"4435",x"4438",x"443B",x"443D",x"4440",x"4442",x"4445",x"4448",x"444A",x"444D",
x"4450",x"4452",x"4455",x"4458",x"445A",x"445D",x"4460",x"4462",x"4465",x"4468",x"446A",x"446D",x"4470",x"4472",x"4475",x"4478",
x"447A",x"447D",x"4480",x"4482",x"4485",x"4488",x"448A",x"448D",x"448F",x"4492",x"4495",x"4497",x"449A",x"449D",x"449F",x"44A2",
x"44A5",x"44A7",x"44AA",x"44AD",x"44AF",x"44B2",x"44B5",x"44B7",x"44BA",x"44BD",x"44BF",x"44C2",x"44C5",x"44C7",x"44CA",x"44CC",
x"44CF",x"44D2",x"44D4",x"44D7",x"44DA",x"44DC",x"44DF",x"44E2",x"44E4",x"44E7",x"44EA",x"44EC",x"44EF",x"44F2",x"44F4",x"44F7",
x"44F9",x"44FC",x"44FF",x"4501",x"4504",x"4507",x"4509",x"450C",x"450F",x"4511",x"4514",x"4517",x"4519",x"451C",x"451F",x"4521",
x"4524",x"4526",x"4529",x"452C",x"452E",x"4531",x"4534",x"4536",x"4539",x"453C",x"453E",x"4541",x"4544",x"4546",x"4549",x"454B",
x"454E",x"4551",x"4553",x"4556",x"4559",x"455B",x"455E",x"4561",x"4563",x"4566",x"4568",x"456B",x"456E",x"4570",x"4573",x"4576",
x"4578",x"457B",x"457E",x"4580",x"4583",x"4586",x"4588",x"458B",x"458D",x"4590",x"4593",x"4595",x"4598",x"459B",x"459D",x"45A0",
x"45A3",x"45A5",x"45A8",x"45AA",x"45AD",x"45B0",x"45B2",x"45B5",x"45B8",x"45BA",x"45BD",x"45BF",x"45C2",x"45C5",x"45C7",x"45CA",
x"45CD",x"45CF",x"45D2",x"45D5",x"45D7",x"45DA",x"45DC",x"45DF",x"45E2",x"45E4",x"45E7",x"45EA",x"45EC",x"45EF",x"45F2",x"45F4",
x"45F7",x"45F9",x"45FC",x"45FF",x"4601",x"4604",x"4607",x"4609",x"460C",x"460E",x"4611",x"4614",x"4616",x"4619",x"461C",x"461E",
x"4621",x"4623",x"4626",x"4629",x"462B",x"462E",x"4631",x"4633",x"4636",x"4638",x"463B",x"463E",x"4640",x"4643",x"4646",x"4648",
x"464B",x"464D",x"4650",x"4653",x"4655",x"4658",x"465B",x"465D",x"4660",x"4662",x"4665",x"4668",x"466A",x"466D",x"4670",x"4672",
x"4675",x"4677",x"467A",x"467D",x"467F",x"4682",x"4685",x"4687",x"468A",x"468C",x"468F",x"4692",x"4694",x"4697",x"469A",x"469C",
x"469F",x"46A1",x"46A4",x"46A7",x"46A9",x"46AC",x"46AF",x"46B1",x"46B4",x"46B6",x"46B9",x"46BC",x"46BE",x"46C1",x"46C3",x"46C6",
x"46C9",x"46CB",x"46CE",x"46D1",x"46D3",x"46D6",x"46D8",x"46DB",x"46DE",x"46E0",x"46E3",x"46E5",x"46E8",x"46EB",x"46ED",x"46F0",
x"46F3",x"46F5",x"46F8",x"46FA",x"46FD",x"4700",x"4702",x"4705",x"4707",x"470A",x"470D",x"470F",x"4712",x"4715",x"4717",x"471A",
x"471C",x"471F",x"4722",x"4724",x"4727",x"4729",x"472C",x"472F",x"4731",x"4734",x"4736",x"4739",x"473C",x"473E",x"4741",x"4744",
x"4746",x"4749",x"474B",x"474E",x"4751",x"4753",x"4756",x"4758",x"475B",x"475E",x"4760",x"4763",x"4765",x"4768",x"476B",x"476D",
x"4770",x"4772",x"4775",x"4778",x"477A",x"477D",x"4780",x"4782",x"4785",x"4787",x"478A",x"478D",x"478F",x"4792",x"4794",x"4797",
x"479A",x"479C",x"479F",x"47A1",x"47A4",x"47A7",x"47A9",x"47AC",x"47AE",x"47B1",x"47B4",x"47B6",x"47B9",x"47BB",x"47BE",x"47C1",
x"47C3",x"47C6",x"47C8",x"47CB",x"47CE",x"47D0",x"47D3",x"47D5",x"47D8",x"47DB",x"47DD",x"47E0",x"47E2",x"47E5",x"47E8",x"47EA",
x"47ED",x"47EF",x"47F2",x"47F5",x"47F7",x"47FA",x"47FC",x"47FF",x"4802",x"4804",x"4807",x"4809",x"480C",x"480F",x"4811",x"4814",
x"4816",x"4819",x"481C",x"481E",x"4821",x"4823",x"4826",x"4829",x"482B",x"482E",x"4830",x"4833",x"4835",x"4838",x"483B",x"483D",
x"4840",x"4842",x"4845",x"4848",x"484A",x"484D",x"484F",x"4852",x"4855",x"4857",x"485A",x"485C",x"485F",x"4862",x"4864",x"4867",
x"4869",x"486C",x"486F",x"4871",x"4874",x"4876",x"4879",x"487B",x"487E",x"4881",x"4883",x"4886",x"4888",x"488B",x"488E",x"4890",
x"4893",x"4895",x"4898",x"489B",x"489D",x"48A0",x"48A2",x"48A5",x"48A7",x"48AA",x"48AD",x"48AF",x"48B2",x"48B4",x"48B7",x"48BA",
x"48BC",x"48BF",x"48C1",x"48C4",x"48C6",x"48C9",x"48CC",x"48CE",x"48D1",x"48D3",x"48D6",x"48D9",x"48DB",x"48DE",x"48E0",x"48E3",
x"48E5",x"48E8",x"48EB",x"48ED",x"48F0",x"48F2",x"48F5",x"48F8",x"48FA",x"48FD",x"48FF",x"4902",x"4904",x"4907",x"490A",x"490C",
x"490F",x"4911",x"4914",x"4917",x"4919",x"491C",x"491E",x"4921",x"4923",x"4926",x"4929",x"492B",x"492E",x"4930",x"4933",x"4935",
x"4938",x"493B",x"493D",x"4940",x"4942",x"4945",x"4947",x"494A",x"494D",x"494F",x"4952",x"4954",x"4957",x"495A",x"495C",x"495F",
x"4961",x"4964",x"4966",x"4969",x"496C",x"496E",x"4971",x"4973",x"4976",x"4978",x"497B",x"497E",x"4980",x"4983",x"4985",x"4988",
x"498A",x"498D",x"4990",x"4992",x"4995",x"4997",x"499A",x"499C",x"499F",x"49A2",x"49A4",x"49A7",x"49A9",x"49AC",x"49AE",x"49B1",
x"49B4",x"49B6",x"49B9",x"49BB",x"49BE",x"49C0",x"49C3",x"49C5",x"49C8",x"49CB",x"49CD",x"49D0",x"49D2",x"49D5",x"49D7",x"49DA",
x"49DD",x"49DF",x"49E2",x"49E4",x"49E7",x"49E9",x"49EC",x"49EF",x"49F1",x"49F4",x"49F6",x"49F9",x"49FB",x"49FE",x"4A00",x"4A03",
x"4A06",x"4A08",x"4A0B",x"4A0D",x"4A10",x"4A12",x"4A15",x"4A18",x"4A1A",x"4A1D",x"4A1F",x"4A22",x"4A24",x"4A27",x"4A29",x"4A2C",
x"4A2F",x"4A31",x"4A34",x"4A36",x"4A39",x"4A3B",x"4A3E",x"4A41",x"4A43",x"4A46",x"4A48",x"4A4B",x"4A4D",x"4A50",x"4A52",x"4A55",
x"4A58",x"4A5A",x"4A5D",x"4A5F",x"4A62",x"4A64",x"4A67",x"4A69",x"4A6C",x"4A6F",x"4A71",x"4A74",x"4A76",x"4A79",x"4A7B",x"4A7E",
x"4A80",x"4A83",x"4A86",x"4A88",x"4A8B",x"4A8D",x"4A90",x"4A92",x"4A95",x"4A97",x"4A9A",x"4A9D",x"4A9F",x"4AA2",x"4AA4",x"4AA7",
x"4AA9",x"4AAC",x"4AAE",x"4AB1",x"4AB3",x"4AB6",x"4AB9",x"4ABB",x"4ABE",x"4AC0",x"4AC3",x"4AC5",x"4AC8",x"4ACA",x"4ACD",x"4AD0",
x"4AD2",x"4AD5",x"4AD7",x"4ADA",x"4ADC",x"4ADF",x"4AE1",x"4AE4",x"4AE6",x"4AE9",x"4AEC",x"4AEE",x"4AF1",x"4AF3",x"4AF6",x"4AF8",
x"4AFB",x"4AFD",x"4B00",x"4B02",x"4B05",x"4B08",x"4B0A",x"4B0D",x"4B0F",x"4B12",x"4B14",x"4B17",x"4B19",x"4B1C",x"4B1E",x"4B21",
x"4B24",x"4B26",x"4B29",x"4B2B",x"4B2E",x"4B30",x"4B33",x"4B35",x"4B38",x"4B3A",x"4B3D",x"4B40",x"4B42",x"4B45",x"4B47",x"4B4A",
x"4B4C",x"4B4F",x"4B51",x"4B54",x"4B56",x"4B59",x"4B5B",x"4B5E",x"4B61",x"4B63",x"4B66",x"4B68",x"4B6B",x"4B6D",x"4B70",x"4B72",
x"4B75",x"4B77",x"4B7A",x"4B7C",x"4B7F",x"4B82",x"4B84",x"4B87",x"4B89",x"4B8C",x"4B8E",x"4B91",x"4B93",x"4B96",x"4B98",x"4B9B",
x"4B9D",x"4BA0",x"4BA2",x"4BA5",x"4BA8",x"4BAA",x"4BAD",x"4BAF",x"4BB2",x"4BB4",x"4BB7",x"4BB9",x"4BBC",x"4BBE",x"4BC1",x"4BC3",
x"4BC6",x"4BC8",x"4BCB",x"4BCE",x"4BD0",x"4BD3",x"4BD5",x"4BD8",x"4BDA",x"4BDD",x"4BDF",x"4BE2",x"4BE4",x"4BE7",x"4BE9",x"4BEC",
x"4BEE",x"4BF1",x"4BF4",x"4BF6",x"4BF9",x"4BFB",x"4BFE",x"4C00",x"4C03",x"4C05",x"4C08",x"4C0A",x"4C0D",x"4C0F",x"4C12",x"4C14",
x"4C17",x"4C19",x"4C1C",x"4C1E",x"4C21",x"4C24",x"4C26",x"4C29",x"4C2B",x"4C2E",x"4C30",x"4C33",x"4C35",x"4C38",x"4C3A",x"4C3D",
x"4C3F",x"4C42",x"4C44",x"4C47",x"4C49",x"4C4C",x"4C4E",x"4C51",x"4C53",x"4C56",x"4C59",x"4C5B",x"4C5E",x"4C60",x"4C63",x"4C65",
x"4C68",x"4C6A",x"4C6D",x"4C6F",x"4C72",x"4C74",x"4C77",x"4C79",x"4C7C",x"4C7E",x"4C81",x"4C83",x"4C86",x"4C88",x"4C8B",x"4C8D",
x"4C90",x"4C92",x"4C95",x"4C97",x"4C9A",x"4C9D",x"4C9F",x"4CA2",x"4CA4",x"4CA7",x"4CA9",x"4CAC",x"4CAE",x"4CB1",x"4CB3",x"4CB6",
x"4CB8",x"4CBB",x"4CBD",x"4CC0",x"4CC2",x"4CC5",x"4CC7",x"4CCA",x"4CCC",x"4CCF",x"4CD1",x"4CD4",x"4CD6",x"4CD9",x"4CDB",x"4CDE",
x"4CE0",x"4CE3",x"4CE5",x"4CE8",x"4CEA",x"4CED",x"4CEF",x"4CF2",x"4CF4",x"4CF7",x"4CFA",x"4CFC",x"4CFF",x"4D01",x"4D04",x"4D06",
x"4D09",x"4D0B",x"4D0E",x"4D10",x"4D13",x"4D15",x"4D18",x"4D1A",x"4D1D",x"4D1F",x"4D22",x"4D24",x"4D27",x"4D29",x"4D2C",x"4D2E",
x"4D31",x"4D33",x"4D36",x"4D38",x"4D3B",x"4D3D",x"4D40",x"4D42",x"4D45",x"4D47",x"4D4A",x"4D4C",x"4D4F",x"4D51",x"4D54",x"4D56",
x"4D59",x"4D5B",x"4D5E",x"4D60",x"4D63",x"4D65",x"4D68",x"4D6A",x"4D6D",x"4D6F",x"4D72",x"4D74",x"4D77",x"4D79",x"4D7C",x"4D7E",
x"4D81",x"4D83",x"4D86",x"4D88",x"4D8B",x"4D8D",x"4D90",x"4D92",x"4D95",x"4D97",x"4D9A",x"4D9C",x"4D9F",x"4DA1",x"4DA4",x"4DA6",
x"4DA9",x"4DAB",x"4DAE",x"4DB0",x"4DB3",x"4DB5",x"4DB8",x"4DBA",x"4DBD",x"4DBF",x"4DC2",x"4DC4",x"4DC7",x"4DC9",x"4DCC",x"4DCE",
x"4DD1",x"4DD3",x"4DD6",x"4DD8",x"4DDB",x"4DDD",x"4DE0",x"4DE2",x"4DE5",x"4DE7",x"4DEA",x"4DEC",x"4DEF",x"4DF1",x"4DF4",x"4DF6",
x"4DF9",x"4DFB",x"4DFE",x"4E00",x"4E03",x"4E05",x"4E08",x"4E0A",x"4E0D",x"4E0F",x"4E11",x"4E14",x"4E16",x"4E19",x"4E1B",x"4E1E",
x"4E20",x"4E23",x"4E25",x"4E28",x"4E2A",x"4E2D",x"4E2F",x"4E32",x"4E34",x"4E37",x"4E39",x"4E3C",x"4E3E",x"4E41",x"4E43",x"4E46",
x"4E48",x"4E4B",x"4E4D",x"4E50",x"4E52",x"4E55",x"4E57",x"4E5A",x"4E5C",x"4E5F",x"4E61",x"4E64",x"4E66",x"4E68",x"4E6B",x"4E6D",
x"4E70",x"4E72",x"4E75",x"4E77",x"4E7A",x"4E7C",x"4E7F",x"4E81",x"4E84",x"4E86",x"4E89",x"4E8B",x"4E8E",x"4E90",x"4E93",x"4E95",
x"4E98",x"4E9A",x"4E9D",x"4E9F",x"4EA2",x"4EA4",x"4EA7",x"4EA9",x"4EAB",x"4EAE",x"4EB0",x"4EB3",x"4EB5",x"4EB8",x"4EBA",x"4EBD",
x"4EBF",x"4EC2",x"4EC4",x"4EC7",x"4EC9",x"4ECC",x"4ECE",x"4ED1",x"4ED3",x"4ED6",x"4ED8",x"4EDB",x"4EDD",x"4EDF",x"4EE2",x"4EE4",
x"4EE7",x"4EE9",x"4EEC",x"4EEE",x"4EF1",x"4EF3",x"4EF6",x"4EF8",x"4EFB",x"4EFD",x"4F00",x"4F02",x"4F05",x"4F07",x"4F0A",x"4F0C",
x"4F0E",x"4F11",x"4F13",x"4F16",x"4F18",x"4F1B",x"4F1D",x"4F20",x"4F22",x"4F25",x"4F27",x"4F2A",x"4F2C",x"4F2F",x"4F31",x"4F33",
x"4F36",x"4F38",x"4F3B",x"4F3D",x"4F40",x"4F42",x"4F45",x"4F47",x"4F4A",x"4F4C",x"4F4F",x"4F51",x"4F54",x"4F56",x"4F58",x"4F5B",
x"4F5D",x"4F60",x"4F62",x"4F65",x"4F67",x"4F6A",x"4F6C",x"4F6F",x"4F71",x"4F74",x"4F76",x"4F79",x"4F7B",x"4F7D",x"4F80",x"4F82",
x"4F85",x"4F87",x"4F8A",x"4F8C",x"4F8F",x"4F91",x"4F94",x"4F96",x"4F99",x"4F9B",x"4F9D",x"4FA0",x"4FA2",x"4FA5",x"4FA7",x"4FAA",
x"4FAC",x"4FAF",x"4FB1",x"4FB4",x"4FB6",x"4FB8",x"4FBB",x"4FBD",x"4FC0",x"4FC2",x"4FC5",x"4FC7",x"4FCA",x"4FCC",x"4FCF",x"4FD1",
x"4FD4",x"4FD6",x"4FD8",x"4FDB",x"4FDD",x"4FE0",x"4FE2",x"4FE5",x"4FE7",x"4FEA",x"4FEC",x"4FEF",x"4FF1",x"4FF3",x"4FF6",x"4FF8",
x"4FFB",x"4FFD",x"5000",x"5002",x"5005",x"5007",x"5009",x"500C",x"500E",x"5011",x"5013",x"5016",x"5018",x"501B",x"501D",x"5020",
x"5022",x"5024",x"5027",x"5029",x"502C",x"502E",x"5031",x"5033",x"5036",x"5038",x"503A",x"503D",x"503F",x"5042",x"5044",x"5047",
x"5049",x"504C",x"504E",x"5050",x"5053",x"5055",x"5058",x"505A",x"505D",x"505F",x"5062",x"5064",x"5067",x"5069",x"506B",x"506E",
x"5070",x"5073",x"5075",x"5078",x"507A",x"507C",x"507F",x"5081",x"5084",x"5086",x"5089",x"508B",x"508E",x"5090",x"5092",x"5095",
x"5097",x"509A",x"509C",x"509F",x"50A1",x"50A4",x"50A6",x"50A8",x"50AB",x"50AD",x"50B0",x"50B2",x"50B5",x"50B7",x"50BA",x"50BC",
x"50BE",x"50C1",x"50C3",x"50C6",x"50C8",x"50CB",x"50CD",x"50CF",x"50D2",x"50D4",x"50D7",x"50D9",x"50DC",x"50DE",x"50E0",x"50E3",
x"50E5",x"50E8",x"50EA",x"50ED",x"50EF",x"50F2",x"50F4",x"50F6",x"50F9",x"50FB",x"50FE",x"5100",x"5103",x"5105",x"5107",x"510A",
x"510C",x"510F",x"5111",x"5114",x"5116",x"5118",x"511B",x"511D",x"5120",x"5122",x"5125",x"5127",x"5129",x"512C",x"512E",x"5131",
x"5133",x"5136",x"5138",x"513A",x"513D",x"513F",x"5142",x"5144",x"5147",x"5149",x"514B",x"514E",x"5150",x"5153",x"5155",x"5158",
x"515A",x"515C",x"515F",x"5161",x"5164",x"5166",x"5169",x"516B",x"516D",x"5170",x"5172",x"5175",x"5177",x"517A",x"517C",x"517E",
x"5181",x"5183",x"5186",x"5188",x"518A",x"518D",x"518F",x"5192",x"5194",x"5197",x"5199",x"519B",x"519E",x"51A0",x"51A3",x"51A5",
x"51A8",x"51AA",x"51AC",x"51AF",x"51B1",x"51B4",x"51B6",x"51B8",x"51BB",x"51BD",x"51C0",x"51C2",x"51C5",x"51C7",x"51C9",x"51CC",
x"51CE",x"51D1",x"51D3",x"51D5",x"51D8",x"51DA",x"51DD",x"51DF",x"51E2",x"51E4",x"51E6",x"51E9",x"51EB",x"51EE",x"51F0",x"51F2",
x"51F5",x"51F7",x"51FA",x"51FC",x"51FE",x"5201",x"5203",x"5206",x"5208",x"520B",x"520D",x"520F",x"5212",x"5214",x"5217",x"5219",
x"521B",x"521E",x"5220",x"5223",x"5225",x"5227",x"522A",x"522C",x"522F",x"5231",x"5233",x"5236",x"5238",x"523B",x"523D",x"5240",
x"5242",x"5244",x"5247",x"5249",x"524C",x"524E",x"5250",x"5253",x"5255",x"5258",x"525A",x"525C",x"525F",x"5261",x"5264",x"5266",
x"5268",x"526B",x"526D",x"5270",x"5272",x"5274",x"5277",x"5279",x"527C",x"527E",x"5280",x"5283",x"5285",x"5288",x"528A",x"528C",
x"528F",x"5291",x"5294",x"5296",x"5298",x"529B",x"529D",x"52A0",x"52A2",x"52A4",x"52A7",x"52A9",x"52AC",x"52AE",x"52B0",x"52B3",
x"52B5",x"52B8",x"52BA",x"52BC",x"52BF",x"52C1",x"52C4",x"52C6",x"52C8",x"52CB",x"52CD",x"52D0",x"52D2",x"52D4",x"52D7",x"52D9",
x"52DC",x"52DE",x"52E0",x"52E3",x"52E5",x"52E8",x"52EA",x"52EC",x"52EF",x"52F1",x"52F4",x"52F6",x"52F8",x"52FB",x"52FD",x"52FF",
x"5302",x"5304",x"5307",x"5309",x"530B",x"530E",x"5310",x"5313",x"5315",x"5317",x"531A",x"531C",x"531F",x"5321",x"5323",x"5326",
x"5328",x"532A",x"532D",x"532F",x"5332",x"5334",x"5336",x"5339",x"533B",x"533E",x"5340",x"5342",x"5345",x"5347",x"534A",x"534C",
x"534E",x"5351",x"5353",x"5355",x"5358",x"535A",x"535D",x"535F",x"5361",x"5364",x"5366",x"5369",x"536B",x"536D",x"5370",x"5372",
x"5374",x"5377",x"5379",x"537C",x"537E",x"5380",x"5383",x"5385",x"5387",x"538A",x"538C",x"538F",x"5391",x"5393",x"5396",x"5398",
x"539B",x"539D",x"539F",x"53A2",x"53A4",x"53A6",x"53A9",x"53AB",x"53AE",x"53B0",x"53B2",x"53B5",x"53B7",x"53B9",x"53BC",x"53BE",
x"53C1",x"53C3",x"53C5",x"53C8",x"53CA",x"53CC",x"53CF",x"53D1",x"53D4",x"53D6",x"53D8",x"53DB",x"53DD",x"53DF",x"53E2",x"53E4",
x"53E7",x"53E9",x"53EB",x"53EE",x"53F0",x"53F2",x"53F5",x"53F7",x"53FA",x"53FC",x"53FE",x"5401",x"5403",x"5405",x"5408",x"540A",
x"540C",x"540F",x"5411",x"5414",x"5416",x"5418",x"541B",x"541D",x"541F",x"5422",x"5424",x"5427",x"5429",x"542B",x"542E",x"5430",
x"5432",x"5435",x"5437",x"5439",x"543C",x"543E",x"5441",x"5443",x"5445",x"5448",x"544A",x"544C",x"544F",x"5451",x"5453",x"5456",
x"5458",x"545B",x"545D",x"545F",x"5462",x"5464",x"5466",x"5469",x"546B",x"546D",x"5470",x"5472",x"5475",x"5477",x"5479",x"547C",
x"547E",x"5480",x"5483",x"5485",x"5487",x"548A",x"548C",x"548E",x"5491",x"5493",x"5496",x"5498",x"549A",x"549D",x"549F",x"54A1",
x"54A4",x"54A6",x"54A8",x"54AB",x"54AD",x"54AF",x"54B2",x"54B4",x"54B7",x"54B9",x"54BB",x"54BE",x"54C0",x"54C2",x"54C5",x"54C7",
x"54C9",x"54CC",x"54CE",x"54D0",x"54D3",x"54D5",x"54D7",x"54DA",x"54DC",x"54DF",x"54E1",x"54E3",x"54E6",x"54E8",x"54EA",x"54ED",
x"54EF",x"54F1",x"54F4",x"54F6",x"54F8",x"54FB",x"54FD",x"54FF",x"5502",x"5504",x"5506",x"5509",x"550B",x"550E",x"5510",x"5512",
x"5515",x"5517",x"5519",x"551C",x"551E",x"5520",x"5523",x"5525",x"5527",x"552A",x"552C",x"552E",x"5531",x"5533",x"5535",x"5538",
x"553A",x"553C",x"553F",x"5541",x"5543",x"5546",x"5548",x"554B",x"554D",x"554F",x"5552",x"5554",x"5556",x"5559",x"555B",x"555D",
x"5560",x"5562",x"5564",x"5567",x"5569",x"556B",x"556E",x"5570",x"5572",x"5575",x"5577",x"5579",x"557C",x"557E",x"5580",x"5583",
x"5585",x"5587",x"558A",x"558C",x"558E",x"5591",x"5593",x"5595",x"5598",x"559A",x"559C",x"559F",x"55A1",x"55A3",x"55A6",x"55A8",
x"55AA",x"55AD",x"55AF",x"55B1",x"55B4",x"55B6",x"55B8",x"55BB",x"55BD",x"55BF",x"55C2",x"55C4",x"55C6",x"55C9",x"55CB",x"55CD",
x"55D0",x"55D2",x"55D4",x"55D7",x"55D9",x"55DB",x"55DE",x"55E0",x"55E2",x"55E5",x"55E7",x"55E9",x"55EC",x"55EE",x"55F0",x"55F3",
x"55F5",x"55F7",x"55FA",x"55FC",x"55FE",x"5601",x"5603",x"5605",x"5608",x"560A",x"560C",x"560F",x"5611",x"5613",x"5616",x"5618",
x"561A",x"561D",x"561F",x"5621",x"5623",x"5626",x"5628",x"562A",x"562D",x"562F",x"5631",x"5634",x"5636",x"5638",x"563B",x"563D",
x"563F",x"5642",x"5644",x"5646",x"5649",x"564B",x"564D",x"5650",x"5652",x"5654",x"5657",x"5659",x"565B",x"565E",x"5660",x"5662",
x"5664",x"5667",x"5669",x"566B",x"566E",x"5670",x"5672",x"5675",x"5677",x"5679",x"567C",x"567E",x"5680",x"5683",x"5685",x"5687",
x"568A",x"568C",x"568E",x"5690",x"5693",x"5695",x"5697",x"569A",x"569C",x"569E",x"56A1",x"56A3",x"56A5",x"56A8",x"56AA",x"56AC",
x"56AF",x"56B1",x"56B3",x"56B5",x"56B8",x"56BA",x"56BC",x"56BF",x"56C1",x"56C3",x"56C6",x"56C8",x"56CA",x"56CD",x"56CF",x"56D1",
x"56D3",x"56D6",x"56D8",x"56DA",x"56DD",x"56DF",x"56E1",x"56E4",x"56E6",x"56E8",x"56EB",x"56ED",x"56EF",x"56F1",x"56F4",x"56F6",
x"56F8",x"56FB",x"56FD",x"56FF",x"5702",x"5704",x"5706",x"5709",x"570B",x"570D",x"570F",x"5712",x"5714",x"5716",x"5719",x"571B",
x"571D",x"5720",x"5722",x"5724",x"5726",x"5729",x"572B",x"572D",x"5730",x"5732",x"5734",x"5737",x"5739",x"573B",x"573D",x"5740",
x"5742",x"5744",x"5747",x"5749",x"574B",x"574E",x"5750",x"5752",x"5754",x"5757",x"5759",x"575B",x"575E",x"5760",x"5762",x"5765",
x"5767",x"5769",x"576B",x"576E",x"5770",x"5772",x"5775",x"5777",x"5779",x"577B",x"577E",x"5780",x"5782",x"5785",x"5787",x"5789",
x"578B",x"578E",x"5790",x"5792",x"5795",x"5797",x"5799",x"579C",x"579E",x"57A0",x"57A2",x"57A5",x"57A7",x"57A9",x"57AC",x"57AE",
x"57B0",x"57B2",x"57B5",x"57B7",x"57B9",x"57BC",x"57BE",x"57C0",x"57C2",x"57C5",x"57C7",x"57C9",x"57CC",x"57CE",x"57D0",x"57D2",
x"57D5",x"57D7",x"57D9",x"57DC",x"57DE",x"57E0",x"57E2",x"57E5",x"57E7",x"57E9",x"57EC",x"57EE",x"57F0",x"57F2",x"57F5",x"57F7",
x"57F9",x"57FC",x"57FE",x"5800",x"5802",x"5805",x"5807",x"5809",x"580C",x"580E",x"5810",x"5812",x"5815",x"5817",x"5819",x"581B",
x"581E",x"5820",x"5822",x"5825",x"5827",x"5829",x"582B",x"582E",x"5830",x"5832",x"5835",x"5837",x"5839",x"583B",x"583E",x"5840",
x"5842",x"5844",x"5847",x"5849",x"584B",x"584E",x"5850",x"5852",x"5854",x"5857",x"5859",x"585B",x"585D",x"5860",x"5862",x"5864",
x"5867",x"5869",x"586B",x"586D",x"5870",x"5872",x"5874",x"5876",x"5879",x"587B",x"587D",x"5880",x"5882",x"5884",x"5886",x"5889",
x"588B",x"588D",x"588F",x"5892",x"5894",x"5896",x"5898",x"589B",x"589D",x"589F",x"58A2",x"58A4",x"58A6",x"58A8",x"58AB",x"58AD",
x"58AF",x"58B1",x"58B4",x"58B6",x"58B8",x"58BA",x"58BD",x"58BF",x"58C1",x"58C4",x"58C6",x"58C8",x"58CA",x"58CD",x"58CF",x"58D1",
x"58D3",x"58D6",x"58D8",x"58DA",x"58DC",x"58DF",x"58E1",x"58E3",x"58E5",x"58E8",x"58EA",x"58EC",x"58EE",x"58F1",x"58F3",x"58F5",
x"58F8",x"58FA",x"58FC",x"58FE",x"5901",x"5903",x"5905",x"5907",x"590A",x"590C",x"590E",x"5910",x"5913",x"5915",x"5917",x"5919",
x"591C",x"591E",x"5920",x"5922",x"5925",x"5927",x"5929",x"592B",x"592E",x"5930",x"5932",x"5934",x"5937",x"5939",x"593B",x"593D",
x"5940",x"5942",x"5944",x"5946",x"5949",x"594B",x"594D",x"594F",x"5952",x"5954",x"5956",x"5958",x"595B",x"595D",x"595F",x"5961",
x"5964",x"5966",x"5968",x"596A",x"596D",x"596F",x"5971",x"5973",x"5976",x"5978",x"597A",x"597C",x"597F",x"5981",x"5983",x"5985",
x"5988",x"598A",x"598C",x"598E",x"5991",x"5993",x"5995",x"5997",x"599A",x"599C",x"599E",x"59A0",x"59A3",x"59A5",x"59A7",x"59A9",
x"59AC",x"59AE",x"59B0",x"59B2",x"59B5",x"59B7",x"59B9",x"59BB",x"59BD",x"59C0",x"59C2",x"59C4",x"59C6",x"59C9",x"59CB",x"59CD",
x"59CF",x"59D2",x"59D4",x"59D6",x"59D8",x"59DB",x"59DD",x"59DF",x"59E1",x"59E4",x"59E6",x"59E8",x"59EA",x"59EC",x"59EF",x"59F1",
x"59F3",x"59F5",x"59F8",x"59FA",x"59FC",x"59FE",x"5A01",x"5A03",x"5A05",x"5A07",x"5A0A",x"5A0C",x"5A0E",x"5A10",x"5A12",x"5A15",
x"5A17",x"5A19",x"5A1B",x"5A1E",x"5A20",x"5A22",x"5A24",x"5A27",x"5A29",x"5A2B",x"5A2D",x"5A2F",x"5A32",x"5A34",x"5A36",x"5A38",
x"5A3B",x"5A3D",x"5A3F",x"5A41",x"5A43",x"5A46",x"5A48",x"5A4A",x"5A4C",x"5A4F",x"5A51",x"5A53",x"5A55",x"5A58",x"5A5A",x"5A5C",
x"5A5E",x"5A60",x"5A63",x"5A65",x"5A67",x"5A69",x"5A6C",x"5A6E",x"5A70",x"5A72",x"5A74",x"5A77",x"5A79",x"5A7B",x"5A7D",x"5A80",
x"5A82",x"5A84",x"5A86",x"5A88",x"5A8B",x"5A8D",x"5A8F",x"5A91",x"5A94",x"5A96",x"5A98",x"5A9A",x"5A9C",x"5A9F",x"5AA1",x"5AA3",
x"5AA5",x"5AA8",x"5AAA",x"5AAC",x"5AAE",x"5AB0",x"5AB3",x"5AB5",x"5AB7",x"5AB9",x"5ABB",x"5ABE",x"5AC0",x"5AC2",x"5AC4",x"5AC7",
x"5AC9",x"5ACB",x"5ACD",x"5ACF",x"5AD2",x"5AD4",x"5AD6",x"5AD8",x"5ADA",x"5ADD",x"5ADF",x"5AE1",x"5AE3",x"5AE6",x"5AE8",x"5AEA",
x"5AEC",x"5AEE",x"5AF1",x"5AF3",x"5AF5",x"5AF7",x"5AF9",x"5AFC",x"5AFE",x"5B00",x"5B02",x"5B04",x"5B07",x"5B09",x"5B0B",x"5B0D",
x"5B0F",x"5B12",x"5B14",x"5B16",x"5B18",x"5B1B",x"5B1D",x"5B1F",x"5B21",x"5B23",x"5B26",x"5B28",x"5B2A",x"5B2C",x"5B2E",x"5B31",
x"5B33",x"5B35",x"5B37",x"5B39",x"5B3C",x"5B3E",x"5B40",x"5B42",x"5B44",x"5B47",x"5B49",x"5B4B",x"5B4D",x"5B4F",x"5B52",x"5B54",
x"5B56",x"5B58",x"5B5A",x"5B5D",x"5B5F",x"5B61",x"5B63",x"5B65",x"5B68",x"5B6A",x"5B6C",x"5B6E",x"5B70",x"5B73",x"5B75",x"5B77",
x"5B79",x"5B7B",x"5B7E",x"5B80",x"5B82",x"5B84",x"5B86",x"5B89",x"5B8B",x"5B8D",x"5B8F",x"5B91",x"5B94",x"5B96",x"5B98",x"5B9A",
x"5B9C",x"5B9F",x"5BA1",x"5BA3",x"5BA5",x"5BA7",x"5BAA",x"5BAC",x"5BAE",x"5BB0",x"5BB2",x"5BB4",x"5BB7",x"5BB9",x"5BBB",x"5BBD",
x"5BBF",x"5BC2",x"5BC4",x"5BC6",x"5BC8",x"5BCA",x"5BCD",x"5BCF",x"5BD1",x"5BD3",x"5BD5",x"5BD8",x"5BDA",x"5BDC",x"5BDE",x"5BE0",
x"5BE2",x"5BE5",x"5BE7",x"5BE9",x"5BEB",x"5BED",x"5BF0",x"5BF2",x"5BF4",x"5BF6",x"5BF8",x"5BFA",x"5BFD",x"5BFF",x"5C01",x"5C03",
x"5C05",x"5C08",x"5C0A",x"5C0C",x"5C0E",x"5C10",x"5C13",x"5C15",x"5C17",x"5C19",x"5C1B",x"5C1D",x"5C20",x"5C22",x"5C24",x"5C26",
x"5C28",x"5C2B",x"5C2D",x"5C2F",x"5C31",x"5C33",x"5C35",x"5C38",x"5C3A",x"5C3C",x"5C3E",x"5C40",x"5C42",x"5C45",x"5C47",x"5C49",
x"5C4B",x"5C4D",x"5C50",x"5C52",x"5C54",x"5C56",x"5C58",x"5C5A",x"5C5D",x"5C5F",x"5C61",x"5C63",x"5C65",x"5C67",x"5C6A",x"5C6C",
x"5C6E",x"5C70",x"5C72",x"5C74",x"5C77",x"5C79",x"5C7B",x"5C7D",x"5C7F",x"5C82",x"5C84",x"5C86",x"5C88",x"5C8A",x"5C8C",x"5C8F",
x"5C91",x"5C93",x"5C95",x"5C97",x"5C99",x"5C9C",x"5C9E",x"5CA0",x"5CA2",x"5CA4",x"5CA6",x"5CA9",x"5CAB",x"5CAD",x"5CAF",x"5CB1",
x"5CB3",x"5CB6",x"5CB8",x"5CBA",x"5CBC",x"5CBE",x"5CC0",x"5CC3",x"5CC5",x"5CC7",x"5CC9",x"5CCB",x"5CCD",x"5CD0",x"5CD2",x"5CD4",
x"5CD6",x"5CD8",x"5CDA",x"5CDD",x"5CDF",x"5CE1",x"5CE3",x"5CE5",x"5CE7",x"5CE9",x"5CEC",x"5CEE",x"5CF0",x"5CF2",x"5CF4",x"5CF6",
x"5CF9",x"5CFB",x"5CFD",x"5CFF",x"5D01",x"5D03",x"5D06",x"5D08",x"5D0A",x"5D0C",x"5D0E",x"5D10",x"5D13",x"5D15",x"5D17",x"5D19",
x"5D1B",x"5D1D",x"5D1F",x"5D22",x"5D24",x"5D26",x"5D28",x"5D2A",x"5D2C",x"5D2F",x"5D31",x"5D33",x"5D35",x"5D37",x"5D39",x"5D3B",
x"5D3E",x"5D40",x"5D42",x"5D44",x"5D46",x"5D48",x"5D4B",x"5D4D",x"5D4F",x"5D51",x"5D53",x"5D55",x"5D57",x"5D5A",x"5D5C",x"5D5E",
x"5D60",x"5D62",x"5D64",x"5D66",x"5D69",x"5D6B",x"5D6D",x"5D6F",x"5D71",x"5D73",x"5D75",x"5D78",x"5D7A",x"5D7C",x"5D7E",x"5D80",
x"5D82",x"5D84",x"5D87",x"5D89",x"5D8B",x"5D8D",x"5D8F",x"5D91",x"5D94",x"5D96",x"5D98",x"5D9A",x"5D9C",x"5D9E",x"5DA0",x"5DA3",
x"5DA5",x"5DA7",x"5DA9",x"5DAB",x"5DAD",x"5DAF",x"5DB1",x"5DB4",x"5DB6",x"5DB8",x"5DBA",x"5DBC",x"5DBE",x"5DC0",x"5DC3",x"5DC5",
x"5DC7",x"5DC9",x"5DCB",x"5DCD",x"5DCF",x"5DD2",x"5DD4",x"5DD6",x"5DD8",x"5DDA",x"5DDC",x"5DDE",x"5DE1",x"5DE3",x"5DE5",x"5DE7",
x"5DE9",x"5DEB",x"5DED",x"5DEF",x"5DF2",x"5DF4",x"5DF6",x"5DF8",x"5DFA",x"5DFC",x"5DFE",x"5E01",x"5E03",x"5E05",x"5E07",x"5E09",
x"5E0B",x"5E0D",x"5E0F",x"5E12",x"5E14",x"5E16",x"5E18",x"5E1A",x"5E1C",x"5E1E",x"5E20",x"5E23",x"5E25",x"5E27",x"5E29",x"5E2B",
x"5E2D",x"5E2F",x"5E32",x"5E34",x"5E36",x"5E38",x"5E3A",x"5E3C",x"5E3E",x"5E40",x"5E43",x"5E45",x"5E47",x"5E49",x"5E4B",x"5E4D",
x"5E4F",x"5E51",x"5E54",x"5E56",x"5E58",x"5E5A",x"5E5C",x"5E5E",x"5E60",x"5E62",x"5E64",x"5E67",x"5E69",x"5E6B",x"5E6D",x"5E6F",
x"5E71",x"5E73",x"5E75",x"5E78",x"5E7A",x"5E7C",x"5E7E",x"5E80",x"5E82",x"5E84",x"5E86",x"5E89",x"5E8B",x"5E8D",x"5E8F",x"5E91",
x"5E93",x"5E95",x"5E97",x"5E99",x"5E9C",x"5E9E",x"5EA0",x"5EA2",x"5EA4",x"5EA6",x"5EA8",x"5EAA",x"5EAD",x"5EAF",x"5EB1",x"5EB3",
x"5EB5",x"5EB7",x"5EB9",x"5EBB",x"5EBD",x"5EC0",x"5EC2",x"5EC4",x"5EC6",x"5EC8",x"5ECA",x"5ECC",x"5ECE",x"5ED0",x"5ED3",x"5ED5",
x"5ED7",x"5ED9",x"5EDB",x"5EDD",x"5EDF",x"5EE1",x"5EE3",x"5EE6",x"5EE8",x"5EEA",x"5EEC",x"5EEE",x"5EF0",x"5EF2",x"5EF4",x"5EF6",
x"5EF8",x"5EFB",x"5EFD",x"5EFF",x"5F01",x"5F03",x"5F05",x"5F07",x"5F09",x"5F0B",x"5F0E",x"5F10",x"5F12",x"5F14",x"5F16",x"5F18",
x"5F1A",x"5F1C",x"5F1E",x"5F20",x"5F23",x"5F25",x"5F27",x"5F29",x"5F2B",x"5F2D",x"5F2F",x"5F31",x"5F33",x"5F35",x"5F38",x"5F3A",
x"5F3C",x"5F3E",x"5F40",x"5F42",x"5F44",x"5F46",x"5F48",x"5F4A",x"5F4D",x"5F4F",x"5F51",x"5F53",x"5F55",x"5F57",x"5F59",x"5F5B",
x"5F5D",x"5F5F",x"5F61",x"5F64",x"5F66",x"5F68",x"5F6A",x"5F6C",x"5F6E",x"5F70",x"5F72",x"5F74",x"5F76",x"5F79",x"5F7B",x"5F7D",
x"5F7F",x"5F81",x"5F83",x"5F85",x"5F87",x"5F89",x"5F8B",x"5F8D",x"5F90",x"5F92",x"5F94",x"5F96",x"5F98",x"5F9A",x"5F9C",x"5F9E",
x"5FA0",x"5FA2",x"5FA4",x"5FA7",x"5FA9",x"5FAB",x"5FAD",x"5FAF",x"5FB1",x"5FB3",x"5FB5",x"5FB7",x"5FB9",x"5FBB",x"5FBD",x"5FC0",
x"5FC2",x"5FC4",x"5FC6",x"5FC8",x"5FCA",x"5FCC",x"5FCE",x"5FD0",x"5FD2",x"5FD4",x"5FD6",x"5FD9",x"5FDB",x"5FDD",x"5FDF",x"5FE1",
x"5FE3",x"5FE5",x"5FE7",x"5FE9",x"5FEB",x"5FED",x"5FEF",x"5FF2",x"5FF4",x"5FF6",x"5FF8",x"5FFA",x"5FFC",x"5FFE",x"6000",x"6002",
x"6004",x"6006",x"6008",x"600A",x"600D",x"600F",x"6011",x"6013",x"6015",x"6017",x"6019",x"601B",x"601D",x"601F",x"6021",x"6023",
x"6025",x"6028",x"602A",x"602C",x"602E",x"6030",x"6032",x"6034",x"6036",x"6038",x"603A",x"603C",x"603E",x"6040",x"6042",x"6045",
x"6047",x"6049",x"604B",x"604D",x"604F",x"6051",x"6053",x"6055",x"6057",x"6059",x"605B",x"605D",x"605F",x"6061",x"6064",x"6066",
x"6068",x"606A",x"606C",x"606E",x"6070",x"6072",x"6074",x"6076",x"6078",x"607A",x"607C",x"607E",x"6080",x"6083",x"6085",x"6087",
x"6089",x"608B",x"608D",x"608F",x"6091",x"6093",x"6095",x"6097",x"6099",x"609B",x"609D",x"609F",x"60A1",x"60A4",x"60A6",x"60A8",
x"60AA",x"60AC",x"60AE",x"60B0",x"60B2",x"60B4",x"60B6",x"60B8",x"60BA",x"60BC",x"60BE",x"60C0",x"60C2",x"60C4",x"60C6",x"60C9",
x"60CB",x"60CD",x"60CF",x"60D1",x"60D3",x"60D5",x"60D7",x"60D9",x"60DB",x"60DD",x"60DF",x"60E1",x"60E3",x"60E5",x"60E7",x"60E9",
x"60EB",x"60EE",x"60F0",x"60F2",x"60F4",x"60F6",x"60F8",x"60FA",x"60FC",x"60FE",x"6100",x"6102",x"6104",x"6106",x"6108",x"610A",
x"610C",x"610E",x"6110",x"6112",x"6114",x"6117",x"6119",x"611B",x"611D",x"611F",x"6121",x"6123",x"6125",x"6127",x"6129",x"612B",
x"612D",x"612F",x"6131",x"6133",x"6135",x"6137",x"6139",x"613B",x"613D",x"613F",x"6141",x"6143",x"6146",x"6148",x"614A",x"614C",
x"614E",x"6150",x"6152",x"6154",x"6156",x"6158",x"615A",x"615C",x"615E",x"6160",x"6162",x"6164",x"6166",x"6168",x"616A",x"616C",
x"616E",x"6170",x"6172",x"6174",x"6176",x"6179",x"617B",x"617D",x"617F",x"6181",x"6183",x"6185",x"6187",x"6189",x"618B",x"618D",
x"618F",x"6191",x"6193",x"6195",x"6197",x"6199",x"619B",x"619D",x"619F",x"61A1",x"61A3",x"61A5",x"61A7",x"61A9",x"61AB",x"61AD",
x"61AF",x"61B1",x"61B3",x"61B5",x"61B8",x"61BA",x"61BC",x"61BE",x"61C0",x"61C2",x"61C4",x"61C6",x"61C8",x"61CA",x"61CC",x"61CE",
x"61D0",x"61D2",x"61D4",x"61D6",x"61D8",x"61DA",x"61DC",x"61DE",x"61E0",x"61E2",x"61E4",x"61E6",x"61E8",x"61EA",x"61EC",x"61EE",
x"61F0",x"61F2",x"61F4",x"61F6",x"61F8",x"61FA",x"61FC",x"61FE",x"6200",x"6202",x"6204",x"6206",x"6208",x"620B",x"620D",x"620F",
x"6211",x"6213",x"6215",x"6217",x"6219",x"621B",x"621D",x"621F",x"6221",x"6223",x"6225",x"6227",x"6229",x"622B",x"622D",x"622F",
x"6231",x"6233",x"6235",x"6237",x"6239",x"623B",x"623D",x"623F",x"6241",x"6243",x"6245",x"6247",x"6249",x"624B",x"624D",x"624F",
x"6251",x"6253",x"6255",x"6257",x"6259",x"625B",x"625D",x"625F",x"6261",x"6263",x"6265",x"6267",x"6269",x"626B",x"626D",x"626F",
x"6271",x"6273",x"6275",x"6277",x"6279",x"627B",x"627D",x"627F",x"6281",x"6283",x"6285",x"6287",x"6289",x"628B",x"628D",x"628F",
x"6291",x"6293",x"6295",x"6297",x"6299",x"629B",x"629D",x"629F",x"62A1",x"62A3",x"62A5",x"62A7",x"62A9",x"62AB",x"62AD",x"62AF",
x"62B1",x"62B3",x"62B5",x"62B7",x"62B9",x"62BB",x"62BD",x"62BF",x"62C1",x"62C3",x"62C5",x"62C7",x"62C9",x"62CB",x"62CD",x"62CF",
x"62D1",x"62D3",x"62D5",x"62D7",x"62D9",x"62DB",x"62DD",x"62DF",x"62E1",x"62E3",x"62E5",x"62E7",x"62E9",x"62EB",x"62ED",x"62EF",
x"62F1",x"62F3",x"62F5",x"62F7",x"62F9",x"62FB",x"62FD",x"62FF",x"6301",x"6303",x"6305",x"6307",x"6309",x"630B",x"630D",x"630F",
x"6311",x"6313",x"6315",x"6317",x"6319",x"631B",x"631D",x"631F",x"6321",x"6323",x"6325",x"6327",x"6329",x"632B",x"632D",x"632F",
x"6331",x"6333",x"6335",x"6337",x"6339",x"633B",x"633D",x"633F",x"6341",x"6343",x"6345",x"6347",x"6349",x"634B",x"634D",x"634F",
x"6351",x"6353",x"6355",x"6357",x"6359",x"635B",x"635D",x"635E",x"6360",x"6362",x"6364",x"6366",x"6368",x"636A",x"636C",x"636E",
x"6370",x"6372",x"6374",x"6376",x"6378",x"637A",x"637C",x"637E",x"6380",x"6382",x"6384",x"6386",x"6388",x"638A",x"638C",x"638E",
x"6390",x"6392",x"6394",x"6396",x"6398",x"639A",x"639C",x"639E",x"63A0",x"63A2",x"63A4",x"63A6",x"63A8",x"63AA",x"63AC",x"63AE",
x"63AF",x"63B1",x"63B3",x"63B5",x"63B7",x"63B9",x"63BB",x"63BD",x"63BF",x"63C1",x"63C3",x"63C5",x"63C7",x"63C9",x"63CB",x"63CD",
x"63CF",x"63D1",x"63D3",x"63D5",x"63D7",x"63D9",x"63DB",x"63DD",x"63DF",x"63E1",x"63E3",x"63E5",x"63E7",x"63E9",x"63EA",x"63EC",
x"63EE",x"63F0",x"63F2",x"63F4",x"63F6",x"63F8",x"63FA",x"63FC",x"63FE",x"6400",x"6402",x"6404",x"6406",x"6408",x"640A",x"640C",
x"640E",x"6410",x"6412",x"6414",x"6416",x"6418",x"641A",x"641C",x"641D",x"641F",x"6421",x"6423",x"6425",x"6427",x"6429",x"642B",
x"642D",x"642F",x"6431",x"6433",x"6435",x"6437",x"6439",x"643B",x"643D",x"643F",x"6441",x"6443",x"6445",x"6447",x"6448",x"644A",
x"644C",x"644E",x"6450",x"6452",x"6454",x"6456",x"6458",x"645A",x"645C",x"645E",x"6460",x"6462",x"6464",x"6466",x"6468",x"646A",
x"646C",x"646E",x"646F",x"6471",x"6473",x"6475",x"6477",x"6479",x"647B",x"647D",x"647F",x"6481",x"6483",x"6485",x"6487",x"6489",
x"648B",x"648D",x"648F",x"6491",x"6492",x"6494",x"6496",x"6498",x"649A",x"649C",x"649E",x"64A0",x"64A2",x"64A4",x"64A6",x"64A8",
x"64AA",x"64AC",x"64AE",x"64B0",x"64B2",x"64B3",x"64B5",x"64B7",x"64B9",x"64BB",x"64BD",x"64BF",x"64C1",x"64C3",x"64C5",x"64C7",
x"64C9",x"64CB",x"64CD",x"64CF",x"64D1",x"64D2",x"64D4",x"64D6",x"64D8",x"64DA",x"64DC",x"64DE",x"64E0",x"64E2",x"64E4",x"64E6",
x"64E8",x"64EA",x"64EC",x"64EE",x"64EF",x"64F1",x"64F3",x"64F5",x"64F7",x"64F9",x"64FB",x"64FD",x"64FF",x"6501",x"6503",x"6505",
x"6507",x"6509",x"650A",x"650C",x"650E",x"6510",x"6512",x"6514",x"6516",x"6518",x"651A",x"651C",x"651E",x"6520",x"6522",x"6524",
x"6525",x"6527",x"6529",x"652B",x"652D",x"652F",x"6531",x"6533",x"6535",x"6537",x"6539",x"653B",x"653D",x"653E",x"6540",x"6542",
x"6544",x"6546",x"6548",x"654A",x"654C",x"654E",x"6550",x"6552",x"6554",x"6556",x"6557",x"6559",x"655B",x"655D",x"655F",x"6561",
x"6563",x"6565",x"6567",x"6569",x"656B",x"656D",x"656E",x"6570",x"6572",x"6574",x"6576",x"6578",x"657A",x"657C",x"657E",x"6580",
x"6582",x"6584",x"6585",x"6587",x"6589",x"658B",x"658D",x"658F",x"6591",x"6593",x"6595",x"6597",x"6599",x"659A",x"659C",x"659E",
x"65A0",x"65A2",x"65A4",x"65A6",x"65A8",x"65AA",x"65AC",x"65AE",x"65AF",x"65B1",x"65B3",x"65B5",x"65B7",x"65B9",x"65BB",x"65BD",
x"65BF",x"65C1",x"65C3",x"65C4",x"65C6",x"65C8",x"65CA",x"65CC",x"65CE",x"65D0",x"65D2",x"65D4",x"65D6",x"65D7",x"65D9",x"65DB",
x"65DD",x"65DF",x"65E1",x"65E3",x"65E5",x"65E7",x"65E9",x"65EA",x"65EC",x"65EE",x"65F0",x"65F2",x"65F4",x"65F6",x"65F8",x"65FA",
x"65FC",x"65FD",x"65FF",x"6601",x"6603",x"6605",x"6607",x"6609",x"660B",x"660D",x"660F",x"6610",x"6612",x"6614",x"6616",x"6618",
x"661A",x"661C",x"661E",x"6620",x"6622",x"6623",x"6625",x"6627",x"6629",x"662B",x"662D",x"662F",x"6631",x"6633",x"6634",x"6636",
x"6638",x"663A",x"663C",x"663E",x"6640",x"6642",x"6644",x"6645",x"6647",x"6649",x"664B",x"664D",x"664F",x"6651",x"6653",x"6655",
x"6656",x"6658",x"665A",x"665C",x"665E",x"6660",x"6662",x"6664",x"6666",x"6667",x"6669",x"666B",x"666D",x"666F",x"6671",x"6673",
x"6675",x"6676",x"6678",x"667A",x"667C",x"667E",x"6680",x"6682",x"6684",x"6686",x"6687",x"6689",x"668B",x"668D",x"668F",x"6691",
x"6693",x"6695",x"6696",x"6698",x"669A",x"669C",x"669E",x"66A0",x"66A2",x"66A4",x"66A5",x"66A7",x"66A9",x"66AB",x"66AD",x"66AF",
x"66B1",x"66B3",x"66B4",x"66B6",x"66B8",x"66BA",x"66BC",x"66BE",x"66C0",x"66C2",x"66C3",x"66C5",x"66C7",x"66C9",x"66CB",x"66CD",
x"66CF",x"66D1",x"66D2",x"66D4",x"66D6",x"66D8",x"66DA",x"66DC",x"66DE",x"66E0",x"66E1",x"66E3",x"66E5",x"66E7",x"66E9",x"66EB",
x"66ED",x"66EE",x"66F0",x"66F2",x"66F4",x"66F6",x"66F8",x"66FA",x"66FC",x"66FD",x"66FF",x"6701",x"6703",x"6705",x"6707",x"6709",
x"670A",x"670C",x"670E",x"6710",x"6712",x"6714",x"6716",x"6718",x"6719",x"671B",x"671D",x"671F",x"6721",x"6723",x"6725",x"6726",
x"6728",x"672A",x"672C",x"672E",x"6730",x"6732",x"6733",x"6735",x"6737",x"6739",x"673B",x"673D",x"673F",x"6740",x"6742",x"6744",
x"6746",x"6748",x"674A",x"674C",x"674D",x"674F",x"6751",x"6753",x"6755",x"6757",x"6759",x"675A",x"675C",x"675E",x"6760",x"6762",
x"6764",x"6765",x"6767",x"6769",x"676B",x"676D",x"676F",x"6771",x"6772",x"6774",x"6776",x"6778",x"677A",x"677C",x"677E",x"677F",
x"6781",x"6783",x"6785",x"6787",x"6789",x"678A",x"678C",x"678E",x"6790",x"6792",x"6794",x"6796",x"6797",x"6799",x"679B",x"679D",
x"679F",x"67A1",x"67A2",x"67A4",x"67A6",x"67A8",x"67AA",x"67AC",x"67AE",x"67AF",x"67B1",x"67B3",x"67B5",x"67B7",x"67B9",x"67BA",
x"67BC",x"67BE",x"67C0",x"67C2",x"67C4",x"67C5",x"67C7",x"67C9",x"67CB",x"67CD",x"67CF",x"67D0",x"67D2",x"67D4",x"67D6",x"67D8",
x"67DA",x"67DC",x"67DD",x"67DF",x"67E1",x"67E3",x"67E5",x"67E7",x"67E8",x"67EA",x"67EC",x"67EE",x"67F0",x"67F2",x"67F3",x"67F5",
x"67F7",x"67F9",x"67FB",x"67FD",x"67FE",x"6800",x"6802",x"6804",x"6806",x"6807",x"6809",x"680B",x"680D",x"680F",x"6811",x"6812",
x"6814",x"6816",x"6818",x"681A",x"681C",x"681D",x"681F",x"6821",x"6823",x"6825",x"6827",x"6828",x"682A",x"682C",x"682E",x"6830",
x"6832",x"6833",x"6835",x"6837",x"6839",x"683B",x"683C",x"683E",x"6840",x"6842",x"6844",x"6846",x"6847",x"6849",x"684B",x"684D",
x"684F",x"6851",x"6852",x"6854",x"6856",x"6858",x"685A",x"685B",x"685D",x"685F",x"6861",x"6863",x"6865",x"6866",x"6868",x"686A",
x"686C",x"686E",x"686F",x"6871",x"6873",x"6875",x"6877",x"6879",x"687A",x"687C",x"687E",x"6880",x"6882",x"6883",x"6885",x"6887",
x"6889",x"688B",x"688C",x"688E",x"6890",x"6892",x"6894",x"6896",x"6897",x"6899",x"689B",x"689D",x"689F",x"68A0",x"68A2",x"68A4",
x"68A6",x"68A8",x"68A9",x"68AB",x"68AD",x"68AF",x"68B1",x"68B2",x"68B4",x"68B6",x"68B8",x"68BA",x"68BB",x"68BD",x"68BF",x"68C1",
x"68C3",x"68C5",x"68C6",x"68C8",x"68CA",x"68CC",x"68CE",x"68CF",x"68D1",x"68D3",x"68D5",x"68D7",x"68D8",x"68DA",x"68DC",x"68DE",
x"68E0",x"68E1",x"68E3",x"68E5",x"68E7",x"68E9",x"68EA",x"68EC",x"68EE",x"68F0",x"68F2",x"68F3",x"68F5",x"68F7",x"68F9",x"68FB",
x"68FC",x"68FE",x"6900",x"6902",x"6904",x"6905",x"6907",x"6909",x"690B",x"690D",x"690E",x"6910",x"6912",x"6914",x"6915",x"6917",
x"6919",x"691B",x"691D",x"691E",x"6920",x"6922",x"6924",x"6926",x"6927",x"6929",x"692B",x"692D",x"692F",x"6930",x"6932",x"6934",
x"6936",x"6938",x"6939",x"693B",x"693D",x"693F",x"6940",x"6942",x"6944",x"6946",x"6948",x"6949",x"694B",x"694D",x"694F",x"6951",
x"6952",x"6954",x"6956",x"6958",x"6959",x"695B",x"695D",x"695F",x"6961",x"6962",x"6964",x"6966",x"6968",x"696A",x"696B",x"696D",
x"696F",x"6971",x"6972",x"6974",x"6976",x"6978",x"697A",x"697B",x"697D",x"697F",x"6981",x"6982",x"6984",x"6986",x"6988",x"698A",
x"698B",x"698D",x"698F",x"6991",x"6992",x"6994",x"6996",x"6998",x"699A",x"699B",x"699D",x"699F",x"69A1",x"69A2",x"69A4",x"69A6",
x"69A8",x"69A9",x"69AB",x"69AD",x"69AF",x"69B1",x"69B2",x"69B4",x"69B6",x"69B8",x"69B9",x"69BB",x"69BD",x"69BF",x"69C1",x"69C2",
x"69C4",x"69C6",x"69C8",x"69C9",x"69CB",x"69CD",x"69CF",x"69D0",x"69D2",x"69D4",x"69D6",x"69D8",x"69D9",x"69DB",x"69DD",x"69DF",
x"69E0",x"69E2",x"69E4",x"69E6",x"69E7",x"69E9",x"69EB",x"69ED",x"69EE",x"69F0",x"69F2",x"69F4",x"69F6",x"69F7",x"69F9",x"69FB",
x"69FD",x"69FE",x"6A00",x"6A02",x"6A04",x"6A05",x"6A07",x"6A09",x"6A0B",x"6A0C",x"6A0E",x"6A10",x"6A12",x"6A13",x"6A15",x"6A17",
x"6A19",x"6A1A",x"6A1C",x"6A1E",x"6A20",x"6A21",x"6A23",x"6A25",x"6A27",x"6A29",x"6A2A",x"6A2C",x"6A2E",x"6A30",x"6A31",x"6A33",
x"6A35",x"6A37",x"6A38",x"6A3A",x"6A3C",x"6A3E",x"6A3F",x"6A41",x"6A43",x"6A45",x"6A46",x"6A48",x"6A4A",x"6A4C",x"6A4D",x"6A4F",
x"6A51",x"6A53",x"6A54",x"6A56",x"6A58",x"6A5A",x"6A5B",x"6A5D",x"6A5F",x"6A61",x"6A62",x"6A64",x"6A66",x"6A68",x"6A69",x"6A6B",
x"6A6D",x"6A6F",x"6A70",x"6A72",x"6A74",x"6A75",x"6A77",x"6A79",x"6A7B",x"6A7C",x"6A7E",x"6A80",x"6A82",x"6A83",x"6A85",x"6A87",
x"6A89",x"6A8A",x"6A8C",x"6A8E",x"6A90",x"6A91",x"6A93",x"6A95",x"6A97",x"6A98",x"6A9A",x"6A9C",x"6A9E",x"6A9F",x"6AA1",x"6AA3",
x"6AA4",x"6AA6",x"6AA8",x"6AAA",x"6AAB",x"6AAD",x"6AAF",x"6AB1",x"6AB2",x"6AB4",x"6AB6",x"6AB8",x"6AB9",x"6ABB",x"6ABD",x"6ABF",
x"6AC0",x"6AC2",x"6AC4",x"6AC5",x"6AC7",x"6AC9",x"6ACB",x"6ACC",x"6ACE",x"6AD0",x"6AD2",x"6AD3",x"6AD5",x"6AD7",x"6AD8",x"6ADA",
x"6ADC",x"6ADE",x"6ADF",x"6AE1",x"6AE3",x"6AE5",x"6AE6",x"6AE8",x"6AEA",x"6AEC",x"6AED",x"6AEF",x"6AF1",x"6AF2",x"6AF4",x"6AF6",
x"6AF8",x"6AF9",x"6AFB",x"6AFD",x"6AFE",x"6B00",x"6B02",x"6B04",x"6B05",x"6B07",x"6B09",x"6B0B",x"6B0C",x"6B0E",x"6B10",x"6B11",
x"6B13",x"6B15",x"6B17",x"6B18",x"6B1A",x"6B1C",x"6B1D",x"6B1F",x"6B21",x"6B23",x"6B24",x"6B26",x"6B28",x"6B2A",x"6B2B",x"6B2D",
x"6B2F",x"6B30",x"6B32",x"6B34",x"6B36",x"6B37",x"6B39",x"6B3B",x"6B3C",x"6B3E",x"6B40",x"6B42",x"6B43",x"6B45",x"6B47",x"6B48",
x"6B4A",x"6B4C",x"6B4E",x"6B4F",x"6B51",x"6B53",x"6B54",x"6B56",x"6B58",x"6B5A",x"6B5B",x"6B5D",x"6B5F",x"6B60",x"6B62",x"6B64",
x"6B65",x"6B67",x"6B69",x"6B6B",x"6B6C",x"6B6E",x"6B70",x"6B71",x"6B73",x"6B75",x"6B77",x"6B78",x"6B7A",x"6B7C",x"6B7D",x"6B7F",
x"6B81",x"6B83",x"6B84",x"6B86",x"6B88",x"6B89",x"6B8B",x"6B8D",x"6B8E",x"6B90",x"6B92",x"6B94",x"6B95",x"6B97",x"6B99",x"6B9A",
x"6B9C",x"6B9E",x"6B9F",x"6BA1",x"6BA3",x"6BA5",x"6BA6",x"6BA8",x"6BAA",x"6BAB",x"6BAD",x"6BAF",x"6BB0",x"6BB2",x"6BB4",x"6BB6",
x"6BB7",x"6BB9",x"6BBB",x"6BBC",x"6BBE",x"6BC0",x"6BC1",x"6BC3",x"6BC5",x"6BC6",x"6BC8",x"6BCA",x"6BCC",x"6BCD",x"6BCF",x"6BD1",
x"6BD2",x"6BD4",x"6BD6",x"6BD7",x"6BD9",x"6BDB",x"6BDD",x"6BDE",x"6BE0",x"6BE2",x"6BE3",x"6BE5",x"6BE7",x"6BE8",x"6BEA",x"6BEC",
x"6BED",x"6BEF",x"6BF1",x"6BF2",x"6BF4",x"6BF6",x"6BF8",x"6BF9",x"6BFB",x"6BFD",x"6BFE",x"6C00",x"6C02",x"6C03",x"6C05",x"6C07",
x"6C08",x"6C0A",x"6C0C",x"6C0D",x"6C0F",x"6C11",x"6C12",x"6C14",x"6C16",x"6C18",x"6C19",x"6C1B",x"6C1D",x"6C1E",x"6C20",x"6C22",
x"6C23",x"6C25",x"6C27",x"6C28",x"6C2A",x"6C2C",x"6C2D",x"6C2F",x"6C31",x"6C32",x"6C34",x"6C36",x"6C37",x"6C39",x"6C3B",x"6C3C",
x"6C3E",x"6C40",x"6C42",x"6C43",x"6C45",x"6C47",x"6C48",x"6C4A",x"6C4C",x"6C4D",x"6C4F",x"6C51",x"6C52",x"6C54",x"6C56",x"6C57",
x"6C59",x"6C5B",x"6C5C",x"6C5E",x"6C60",x"6C61",x"6C63",x"6C65",x"6C66",x"6C68",x"6C6A",x"6C6B",x"6C6D",x"6C6F",x"6C70",x"6C72",
x"6C74",x"6C75",x"6C77",x"6C79",x"6C7A",x"6C7C",x"6C7E",x"6C7F",x"6C81",x"6C83",x"6C84",x"6C86",x"6C88",x"6C89",x"6C8B",x"6C8D",
x"6C8E",x"6C90",x"6C92",x"6C93",x"6C95",x"6C97",x"6C98",x"6C9A",x"6C9C",x"6C9D",x"6C9F",x"6CA1",x"6CA2",x"6CA4",x"6CA6",x"6CA7",
x"6CA9",x"6CAB",x"6CAC",x"6CAE",x"6CB0",x"6CB1",x"6CB3",x"6CB5",x"6CB6",x"6CB8",x"6CBA",x"6CBB",x"6CBD",x"6CBF",x"6CC0",x"6CC2",
x"6CC3",x"6CC5",x"6CC7",x"6CC8",x"6CCA",x"6CCC",x"6CCD",x"6CCF",x"6CD1",x"6CD2",x"6CD4",x"6CD6",x"6CD7",x"6CD9",x"6CDB",x"6CDC",
x"6CDE",x"6CE0",x"6CE1",x"6CE3",x"6CE5",x"6CE6",x"6CE8",x"6CEA",x"6CEB",x"6CED",x"6CEE",x"6CF0",x"6CF2",x"6CF3",x"6CF5",x"6CF7",
x"6CF8",x"6CFA",x"6CFC",x"6CFD",x"6CFF",x"6D01",x"6D02",x"6D04",x"6D06",x"6D07",x"6D09",x"6D0A",x"6D0C",x"6D0E",x"6D0F",x"6D11",
x"6D13",x"6D14",x"6D16",x"6D18",x"6D19",x"6D1B",x"6D1D",x"6D1E",x"6D20",x"6D21",x"6D23",x"6D25",x"6D26",x"6D28",x"6D2A",x"6D2B",
x"6D2D",x"6D2F",x"6D30",x"6D32",x"6D34",x"6D35",x"6D37",x"6D38",x"6D3A",x"6D3C",x"6D3D",x"6D3F",x"6D41",x"6D42",x"6D44",x"6D46",
x"6D47",x"6D49",x"6D4A",x"6D4C",x"6D4E",x"6D4F",x"6D51",x"6D53",x"6D54",x"6D56",x"6D58",x"6D59",x"6D5B",x"6D5C",x"6D5E",x"6D60",
x"6D61",x"6D63",x"6D65",x"6D66",x"6D68",x"6D69",x"6D6B",x"6D6D",x"6D6E",x"6D70",x"6D72",x"6D73",x"6D75",x"6D76",x"6D78",x"6D7A",
x"6D7B",x"6D7D",x"6D7F",x"6D80",x"6D82",x"6D84",x"6D85",x"6D87",x"6D88",x"6D8A",x"6D8C",x"6D8D",x"6D8F",x"6D91",x"6D92",x"6D94",
x"6D95",x"6D97",x"6D99",x"6D9A",x"6D9C",x"6D9D",x"6D9F",x"6DA1",x"6DA2",x"6DA4",x"6DA6",x"6DA7",x"6DA9",x"6DAA",x"6DAC",x"6DAE",
x"6DAF",x"6DB1",x"6DB3",x"6DB4",x"6DB6",x"6DB7",x"6DB9",x"6DBB",x"6DBC",x"6DBE",x"6DBF",x"6DC1",x"6DC3",x"6DC4",x"6DC6",x"6DC8",
x"6DC9",x"6DCB",x"6DCC",x"6DCE",x"6DD0",x"6DD1",x"6DD3",x"6DD4",x"6DD6",x"6DD8",x"6DD9",x"6DDB",x"6DDD",x"6DDE",x"6DE0",x"6DE1",
x"6DE3",x"6DE5",x"6DE6",x"6DE8",x"6DE9",x"6DEB",x"6DED",x"6DEE",x"6DF0",x"6DF1",x"6DF3",x"6DF5",x"6DF6",x"6DF8",x"6DFA",x"6DFB",
x"6DFD",x"6DFE",x"6E00",x"6E02",x"6E03",x"6E05",x"6E06",x"6E08",x"6E0A",x"6E0B",x"6E0D",x"6E0E",x"6E10",x"6E12",x"6E13",x"6E15",
x"6E16",x"6E18",x"6E1A",x"6E1B",x"6E1D",x"6E1E",x"6E20",x"6E22",x"6E23",x"6E25",x"6E26",x"6E28",x"6E2A",x"6E2B",x"6E2D",x"6E2E",
x"6E30",x"6E32",x"6E33",x"6E35",x"6E36",x"6E38",x"6E3A",x"6E3B",x"6E3D",x"6E3E",x"6E40",x"6E42",x"6E43",x"6E45",x"6E46",x"6E48",
x"6E4A",x"6E4B",x"6E4D",x"6E4E",x"6E50",x"6E52",x"6E53",x"6E55",x"6E56",x"6E58",x"6E59",x"6E5B",x"6E5D",x"6E5E",x"6E60",x"6E61",
x"6E63",x"6E65",x"6E66",x"6E68",x"6E69",x"6E6B",x"6E6D",x"6E6E",x"6E70",x"6E71",x"6E73",x"6E75",x"6E76",x"6E78",x"6E79",x"6E7B",
x"6E7C",x"6E7E",x"6E80",x"6E81",x"6E83",x"6E84",x"6E86",x"6E88",x"6E89",x"6E8B",x"6E8C",x"6E8E",x"6E8F",x"6E91",x"6E93",x"6E94",
x"6E96",x"6E97",x"6E99",x"6E9B",x"6E9C",x"6E9E",x"6E9F",x"6EA1",x"6EA2",x"6EA4",x"6EA6",x"6EA7",x"6EA9",x"6EAA",x"6EAC",x"6EAD",
x"6EAF",x"6EB1",x"6EB2",x"6EB4",x"6EB5",x"6EB7",x"6EB9",x"6EBA",x"6EBC",x"6EBD",x"6EBF",x"6EC0",x"6EC2",x"6EC4",x"6EC5",x"6EC7",
x"6EC8",x"6ECA",x"6ECB",x"6ECD",x"6ECF",x"6ED0",x"6ED2",x"6ED3",x"6ED5",x"6ED6",x"6ED8",x"6EDA",x"6EDB",x"6EDD",x"6EDE",x"6EE0",
x"6EE1",x"6EE3",x"6EE5",x"6EE6",x"6EE8",x"6EE9",x"6EEB",x"6EEC",x"6EEE",x"6EF0",x"6EF1",x"6EF3",x"6EF4",x"6EF6",x"6EF7",x"6EF9",
x"6EFB",x"6EFC",x"6EFE",x"6EFF",x"6F01",x"6F02",x"6F04",x"6F05",x"6F07",x"6F09",x"6F0A",x"6F0C",x"6F0D",x"6F0F",x"6F10",x"6F12",
x"6F14",x"6F15",x"6F17",x"6F18",x"6F1A",x"6F1B",x"6F1D",x"6F1E",x"6F20",x"6F22",x"6F23",x"6F25",x"6F26",x"6F28",x"6F29",x"6F2B",
x"6F2C",x"6F2E",x"6F30",x"6F31",x"6F33",x"6F34",x"6F36",x"6F37",x"6F39",x"6F3A",x"6F3C",x"6F3E",x"6F3F",x"6F41",x"6F42",x"6F44",
x"6F45",x"6F47",x"6F48",x"6F4A",x"6F4C",x"6F4D",x"6F4F",x"6F50",x"6F52",x"6F53",x"6F55",x"6F56",x"6F58",x"6F59",x"6F5B",x"6F5D",
x"6F5E",x"6F60",x"6F61",x"6F63",x"6F64",x"6F66",x"6F67",x"6F69",x"6F6B",x"6F6C",x"6F6E",x"6F6F",x"6F71",x"6F72",x"6F74",x"6F75",
x"6F77",x"6F78",x"6F7A",x"6F7C",x"6F7D",x"6F7F",x"6F80",x"6F82",x"6F83",x"6F85",x"6F86",x"6F88",x"6F89",x"6F8B",x"6F8C",x"6F8E",
x"6F90",x"6F91",x"6F93",x"6F94",x"6F96",x"6F97",x"6F99",x"6F9A",x"6F9C",x"6F9D",x"6F9F",x"6FA0",x"6FA2",x"6FA4",x"6FA5",x"6FA7",
x"6FA8",x"6FAA",x"6FAB",x"6FAD",x"6FAE",x"6FB0",x"6FB1",x"6FB3",x"6FB4",x"6FB6",x"6FB8",x"6FB9",x"6FBB",x"6FBC",x"6FBE",x"6FBF",
x"6FC1",x"6FC2",x"6FC4",x"6FC5",x"6FC7",x"6FC8",x"6FCA",x"6FCB",x"6FCD",x"6FCE",x"6FD0",x"6FD2",x"6FD3",x"6FD5",x"6FD6",x"6FD8",
x"6FD9",x"6FDB",x"6FDC",x"6FDE",x"6FDF",x"6FE1",x"6FE2",x"6FE4",x"6FE5",x"6FE7",x"6FE8",x"6FEA",x"6FEB",x"6FED",x"6FEF",x"6FF0",
x"6FF2",x"6FF3",x"6FF5",x"6FF6",x"6FF8",x"6FF9",x"6FFB",x"6FFC",x"6FFE",x"6FFF",x"7001",x"7002",x"7004",x"7005",x"7007",x"7008",
x"700A",x"700B",x"700D",x"700E",x"7010",x"7012",x"7013",x"7015",x"7016",x"7018",x"7019",x"701B",x"701C",x"701E",x"701F",x"7021",
x"7022",x"7024",x"7025",x"7027",x"7028",x"702A",x"702B",x"702D",x"702E",x"7030",x"7031",x"7033",x"7034",x"7036",x"7037",x"7039",
x"703A",x"703C",x"703D",x"703F",x"7040",x"7042",x"7043",x"7045",x"7046",x"7048",x"7049",x"704B",x"704C",x"704E",x"7050",x"7051",
x"7053",x"7054",x"7056",x"7057",x"7059",x"705A",x"705C",x"705D",x"705F",x"7060",x"7062",x"7063",x"7065",x"7066",x"7068",x"7069",
x"706B",x"706C",x"706E",x"706F",x"7071",x"7072",x"7074",x"7075",x"7077",x"7078",x"707A",x"707B",x"707D",x"707E",x"7080",x"7081",
x"7083",x"7084",x"7086",x"7087",x"7089",x"708A",x"708C",x"708D",x"708F",x"7090",x"7092",x"7093",x"7095",x"7096",x"7098",x"7099",
x"709B",x"709C",x"709E",x"709F",x"70A0",x"70A2",x"70A3",x"70A5",x"70A6",x"70A8",x"70A9",x"70AB",x"70AC",x"70AE",x"70AF",x"70B1",
x"70B2",x"70B4",x"70B5",x"70B7",x"70B8",x"70BA",x"70BB",x"70BD",x"70BE",x"70C0",x"70C1",x"70C3",x"70C4",x"70C6",x"70C7",x"70C9",
x"70CA",x"70CC",x"70CD",x"70CF",x"70D0",x"70D2",x"70D3",x"70D5",x"70D6",x"70D8",x"70D9",x"70DB",x"70DC",x"70DD",x"70DF",x"70E0",
x"70E2",x"70E3",x"70E5",x"70E6",x"70E8",x"70E9",x"70EB",x"70EC",x"70EE",x"70EF",x"70F1",x"70F2",x"70F4",x"70F5",x"70F7",x"70F8",
x"70FA",x"70FB",x"70FD",x"70FE",x"70FF",x"7101",x"7102",x"7104",x"7105",x"7107",x"7108",x"710A",x"710B",x"710D",x"710E",x"7110",
x"7111",x"7113",x"7114",x"7116",x"7117",x"7119",x"711A",x"711B",x"711D",x"711E",x"7120",x"7121",x"7123",x"7124",x"7126",x"7127",
x"7129",x"712A",x"712C",x"712D",x"712F",x"7130",x"7131",x"7133",x"7134",x"7136",x"7137",x"7139",x"713A",x"713C",x"713D",x"713F",
x"7140",x"7142",x"7143",x"7145",x"7146",x"7147",x"7149",x"714A",x"714C",x"714D",x"714F",x"7150",x"7152",x"7153",x"7155",x"7156",
x"7158",x"7159",x"715A",x"715C",x"715D",x"715F",x"7160",x"7162",x"7163",x"7165",x"7166",x"7168",x"7169",x"716A",x"716C",x"716D",
x"716F",x"7170",x"7172",x"7173",x"7175",x"7176",x"7178",x"7179",x"717A",x"717C",x"717D",x"717F",x"7180",x"7182",x"7183",x"7185",
x"7186",x"7188",x"7189",x"718A",x"718C",x"718D",x"718F",x"7190",x"7192",x"7193",x"7195",x"7196",x"7197",x"7199",x"719A",x"719C",
x"719D",x"719F",x"71A0",x"71A2",x"71A3",x"71A5",x"71A6",x"71A7",x"71A9",x"71AA",x"71AC",x"71AD",x"71AF",x"71B0",x"71B2",x"71B3",
x"71B4",x"71B6",x"71B7",x"71B9",x"71BA",x"71BC",x"71BD",x"71BE",x"71C0",x"71C1",x"71C3",x"71C4",x"71C6",x"71C7",x"71C9",x"71CA",
x"71CB",x"71CD",x"71CE",x"71D0",x"71D1",x"71D3",x"71D4",x"71D6",x"71D7",x"71D8",x"71DA",x"71DB",x"71DD",x"71DE",x"71E0",x"71E1",
x"71E2",x"71E4",x"71E5",x"71E7",x"71E8",x"71EA",x"71EB",x"71EC",x"71EE",x"71EF",x"71F1",x"71F2",x"71F4",x"71F5",x"71F6",x"71F8",
x"71F9",x"71FB",x"71FC",x"71FE",x"71FF",x"7200",x"7202",x"7203",x"7205",x"7206",x"7208",x"7209",x"720A",x"720C",x"720D",x"720F",
x"7210",x"7212",x"7213",x"7214",x"7216",x"7217",x"7219",x"721A",x"721C",x"721D",x"721E",x"7220",x"7221",x"7223",x"7224",x"7226",
x"7227",x"7228",x"722A",x"722B",x"722D",x"722E",x"722F",x"7231",x"7232",x"7234",x"7235",x"7237",x"7238",x"7239",x"723B",x"723C",
x"723E",x"723F",x"7240",x"7242",x"7243",x"7245",x"7246",x"7248",x"7249",x"724A",x"724C",x"724D",x"724F",x"7250",x"7251",x"7253",
x"7254",x"7256",x"7257",x"7259",x"725A",x"725B",x"725D",x"725E",x"7260",x"7261",x"7262",x"7264",x"7265",x"7267",x"7268",x"7269",
x"726B",x"726C",x"726E",x"726F",x"7270",x"7272",x"7273",x"7275",x"7276",x"7278",x"7279",x"727A",x"727C",x"727D",x"727F",x"7280",
x"7281",x"7283",x"7284",x"7286",x"7287",x"7288",x"728A",x"728B",x"728D",x"728E",x"728F",x"7291",x"7292",x"7294",x"7295",x"7296",
x"7298",x"7299",x"729B",x"729C",x"729D",x"729F",x"72A0",x"72A2",x"72A3",x"72A4",x"72A6",x"72A7",x"72A9",x"72AA",x"72AB",x"72AD",
x"72AE",x"72B0",x"72B1",x"72B2",x"72B4",x"72B5",x"72B6",x"72B8",x"72B9",x"72BB",x"72BC",x"72BD",x"72BF",x"72C0",x"72C2",x"72C3",
x"72C4",x"72C6",x"72C7",x"72C9",x"72CA",x"72CB",x"72CD",x"72CE",x"72D0",x"72D1",x"72D2",x"72D4",x"72D5",x"72D6",x"72D8",x"72D9",
x"72DB",x"72DC",x"72DD",x"72DF",x"72E0",x"72E2",x"72E3",x"72E4",x"72E6",x"72E7",x"72E8",x"72EA",x"72EB",x"72ED",x"72EE",x"72EF",
x"72F1",x"72F2",x"72F4",x"72F5",x"72F6",x"72F8",x"72F9",x"72FA",x"72FC",x"72FD",x"72FF",x"7300",x"7301",x"7303",x"7304",x"7305",
x"7307",x"7308",x"730A",x"730B",x"730C",x"730E",x"730F",x"7311",x"7312",x"7313",x"7315",x"7316",x"7317",x"7319",x"731A",x"731C",
x"731D",x"731E",x"7320",x"7321",x"7322",x"7324",x"7325",x"7326",x"7328",x"7329",x"732B",x"732C",x"732D",x"732F",x"7330",x"7331",
x"7333",x"7334",x"7336",x"7337",x"7338",x"733A",x"733B",x"733C",x"733E",x"733F",x"7340",x"7342",x"7343",x"7345",x"7346",x"7347",
x"7349",x"734A",x"734B",x"734D",x"734E",x"7350",x"7351",x"7352",x"7354",x"7355",x"7356",x"7358",x"7359",x"735A",x"735C",x"735D",
x"735E",x"7360",x"7361",x"7363",x"7364",x"7365",x"7367",x"7368",x"7369",x"736B",x"736C",x"736D",x"736F",x"7370",x"7372",x"7373",
x"7374",x"7376",x"7377",x"7378",x"737A",x"737B",x"737C",x"737E",x"737F",x"7380",x"7382",x"7383",x"7384",x"7386",x"7387",x"7389",
x"738A",x"738B",x"738D",x"738E",x"738F",x"7391",x"7392",x"7393",x"7395",x"7396",x"7397",x"7399",x"739A",x"739B",x"739D",x"739E",
x"739F",x"73A1",x"73A2",x"73A4",x"73A5",x"73A6",x"73A8",x"73A9",x"73AA",x"73AC",x"73AD",x"73AE",x"73B0",x"73B1",x"73B2",x"73B4",
x"73B5",x"73B6",x"73B8",x"73B9",x"73BA",x"73BC",x"73BD",x"73BE",x"73C0",x"73C1",x"73C2",x"73C4",x"73C5",x"73C6",x"73C8",x"73C9",
x"73CA",x"73CC",x"73CD",x"73CE",x"73D0",x"73D1",x"73D3",x"73D4",x"73D5",x"73D7",x"73D8",x"73D9",x"73DB",x"73DC",x"73DD",x"73DF",
x"73E0",x"73E1",x"73E3",x"73E4",x"73E5",x"73E7",x"73E8",x"73E9",x"73EB",x"73EC",x"73ED",x"73EF",x"73F0",x"73F1",x"73F3",x"73F4",
x"73F5",x"73F7",x"73F8",x"73F9",x"73FA",x"73FC",x"73FD",x"73FE",x"7400",x"7401",x"7402",x"7404",x"7405",x"7406",x"7408",x"7409",
x"740A",x"740C",x"740D",x"740E",x"7410",x"7411",x"7412",x"7414",x"7415",x"7416",x"7418",x"7419",x"741A",x"741C",x"741D",x"741E",
x"7420",x"7421",x"7422",x"7424",x"7425",x"7426",x"7428",x"7429",x"742A",x"742B",x"742D",x"742E",x"742F",x"7431",x"7432",x"7433",
x"7435",x"7436",x"7437",x"7439",x"743A",x"743B",x"743D",x"743E",x"743F",x"7441",x"7442",x"7443",x"7444",x"7446",x"7447",x"7448",
x"744A",x"744B",x"744C",x"744E",x"744F",x"7450",x"7452",x"7453",x"7454",x"7456",x"7457",x"7458",x"7459",x"745B",x"745C",x"745D",
x"745F",x"7460",x"7461",x"7463",x"7464",x"7465",x"7467",x"7468",x"7469",x"746A",x"746C",x"746D",x"746E",x"7470",x"7471",x"7472",
x"7474",x"7475",x"7476",x"7478",x"7479",x"747A",x"747B",x"747D",x"747E",x"747F",x"7481",x"7482",x"7483",x"7485",x"7486",x"7487",
x"7488",x"748A",x"748B",x"748C",x"748E",x"748F",x"7490",x"7492",x"7493",x"7494",x"7495",x"7497",x"7498",x"7499",x"749B",x"749C",
x"749D",x"749E",x"74A0",x"74A1",x"74A2",x"74A4",x"74A5",x"74A6",x"74A8",x"74A9",x"74AA",x"74AB",x"74AD",x"74AE",x"74AF",x"74B1",
x"74B2",x"74B3",x"74B4",x"74B6",x"74B7",x"74B8",x"74BA",x"74BB",x"74BC",x"74BD",x"74BF",x"74C0",x"74C1",x"74C3",x"74C4",x"74C5",
x"74C6",x"74C8",x"74C9",x"74CA",x"74CC",x"74CD",x"74CE",x"74CF",x"74D1",x"74D2",x"74D3",x"74D5",x"74D6",x"74D7",x"74D8",x"74DA",
x"74DB",x"74DC",x"74DE",x"74DF",x"74E0",x"74E1",x"74E3",x"74E4",x"74E5",x"74E7",x"74E8",x"74E9",x"74EA",x"74EC",x"74ED",x"74EE",
x"74F0",x"74F1",x"74F2",x"74F3",x"74F5",x"74F6",x"74F7",x"74F8",x"74FA",x"74FB",x"74FC",x"74FE",x"74FF",x"7500",x"7501",x"7503",
x"7504",x"7505",x"7506",x"7508",x"7509",x"750A",x"750C",x"750D",x"750E",x"750F",x"7511",x"7512",x"7513",x"7514",x"7516",x"7517",
x"7518",x"751A",x"751B",x"751C",x"751D",x"751F",x"7520",x"7521",x"7522",x"7524",x"7525",x"7526",x"7527",x"7529",x"752A",x"752B",
x"752D",x"752E",x"752F",x"7530",x"7532",x"7533",x"7534",x"7535",x"7537",x"7538",x"7539",x"753A",x"753C",x"753D",x"753E",x"753F",
x"7541",x"7542",x"7543",x"7544",x"7546",x"7547",x"7548",x"754A",x"754B",x"754C",x"754D",x"754F",x"7550",x"7551",x"7552",x"7554",
x"7555",x"7556",x"7557",x"7559",x"755A",x"755B",x"755C",x"755E",x"755F",x"7560",x"7561",x"7563",x"7564",x"7565",x"7566",x"7568",
x"7569",x"756A",x"756B",x"756D",x"756E",x"756F",x"7570",x"7572",x"7573",x"7574",x"7575",x"7577",x"7578",x"7579",x"757A",x"757C",
x"757D",x"757E",x"757F",x"7581",x"7582",x"7583",x"7584",x"7586",x"7587",x"7588",x"7589",x"758B",x"758C",x"758D",x"758E",x"7590",
x"7591",x"7592",x"7593",x"7594",x"7596",x"7597",x"7598",x"7599",x"759B",x"759C",x"759D",x"759E",x"75A0",x"75A1",x"75A2",x"75A3",
x"75A5",x"75A6",x"75A7",x"75A8",x"75AA",x"75AB",x"75AC",x"75AD",x"75AE",x"75B0",x"75B1",x"75B2",x"75B3",x"75B5",x"75B6",x"75B7",
x"75B8",x"75BA",x"75BB",x"75BC",x"75BD",x"75BF",x"75C0",x"75C1",x"75C2",x"75C3",x"75C5",x"75C6",x"75C7",x"75C8",x"75CA",x"75CB",
x"75CC",x"75CD",x"75CF",x"75D0",x"75D1",x"75D2",x"75D3",x"75D5",x"75D6",x"75D7",x"75D8",x"75DA",x"75DB",x"75DC",x"75DD",x"75DE",
x"75E0",x"75E1",x"75E2",x"75E3",x"75E5",x"75E6",x"75E7",x"75E8",x"75E9",x"75EB",x"75EC",x"75ED",x"75EE",x"75F0",x"75F1",x"75F2",
x"75F3",x"75F4",x"75F6",x"75F7",x"75F8",x"75F9",x"75FB",x"75FC",x"75FD",x"75FE",x"75FF",x"7601",x"7602",x"7603",x"7604",x"7606",
x"7607",x"7608",x"7609",x"760A",x"760C",x"760D",x"760E",x"760F",x"7610",x"7612",x"7613",x"7614",x"7615",x"7617",x"7618",x"7619",
x"761A",x"761B",x"761D",x"761E",x"761F",x"7620",x"7621",x"7623",x"7624",x"7625",x"7626",x"7627",x"7629",x"762A",x"762B",x"762C",
x"762D",x"762F",x"7630",x"7631",x"7632",x"7634",x"7635",x"7636",x"7637",x"7638",x"763A",x"763B",x"763C",x"763D",x"763E",x"7640",
x"7641",x"7642",x"7643",x"7644",x"7646",x"7647",x"7648",x"7649",x"764A",x"764C",x"764D",x"764E",x"764F",x"7650",x"7652",x"7653",
x"7654",x"7655",x"7656",x"7658",x"7659",x"765A",x"765B",x"765C",x"765E",x"765F",x"7660",x"7661",x"7662",x"7664",x"7665",x"7666",
x"7667",x"7668",x"7669",x"766B",x"766C",x"766D",x"766E",x"766F",x"7671",x"7672",x"7673",x"7674",x"7675",x"7677",x"7678",x"7679",
x"767A",x"767B",x"767D",x"767E",x"767F",x"7680",x"7681",x"7682",x"7684",x"7685",x"7686",x"7687",x"7688",x"768A",x"768B",x"768C",
x"768D",x"768E",x"768F",x"7691",x"7692",x"7693",x"7694",x"7695",x"7697",x"7698",x"7699",x"769A",x"769B",x"769D",x"769E",x"769F",
x"76A0",x"76A1",x"76A2",x"76A4",x"76A5",x"76A6",x"76A7",x"76A8",x"76A9",x"76AB",x"76AC",x"76AD",x"76AE",x"76AF",x"76B1",x"76B2",
x"76B3",x"76B4",x"76B5",x"76B6",x"76B8",x"76B9",x"76BA",x"76BB",x"76BC",x"76BD",x"76BF",x"76C0",x"76C1",x"76C2",x"76C3",x"76C4",
x"76C6",x"76C7",x"76C8",x"76C9",x"76CA",x"76CC",x"76CD",x"76CE",x"76CF",x"76D0",x"76D1",x"76D3",x"76D4",x"76D5",x"76D6",x"76D7",
x"76D8",x"76DA",x"76DB",x"76DC",x"76DD",x"76DE",x"76DF",x"76E1",x"76E2",x"76E3",x"76E4",x"76E5",x"76E6",x"76E7",x"76E9",x"76EA",
x"76EB",x"76EC",x"76ED",x"76EE",x"76F0",x"76F1",x"76F2",x"76F3",x"76F4",x"76F5",x"76F7",x"76F8",x"76F9",x"76FA",x"76FB",x"76FC",
x"76FE",x"76FF",x"7700",x"7701",x"7702",x"7703",x"7704",x"7706",x"7707",x"7708",x"7709",x"770A",x"770B",x"770D",x"770E",x"770F",
x"7710",x"7711",x"7712",x"7713",x"7715",x"7716",x"7717",x"7718",x"7719",x"771A",x"771C",x"771D",x"771E",x"771F",x"7720",x"7721",
x"7722",x"7724",x"7725",x"7726",x"7727",x"7728",x"7729",x"772A",x"772C",x"772D",x"772E",x"772F",x"7730",x"7731",x"7732",x"7734",
x"7735",x"7736",x"7737",x"7738",x"7739",x"773A",x"773C",x"773D",x"773E",x"773F",x"7740",x"7741",x"7742",x"7744",x"7745",x"7746",
x"7747",x"7748",x"7749",x"774A",x"774C",x"774D",x"774E",x"774F",x"7750",x"7751",x"7752",x"7754",x"7755",x"7756",x"7757",x"7758",
x"7759",x"775A",x"775C",x"775D",x"775E",x"775F",x"7760",x"7761",x"7762",x"7763",x"7765",x"7766",x"7767",x"7768",x"7769",x"776A",
x"776B",x"776D",x"776E",x"776F",x"7770",x"7771",x"7772",x"7773",x"7774",x"7776",x"7777",x"7778",x"7779",x"777A",x"777B",x"777C",
x"777D",x"777F",x"7780",x"7781",x"7782",x"7783",x"7784",x"7785",x"7786",x"7788",x"7789",x"778A",x"778B",x"778C",x"778D",x"778E",
x"778F",x"7791",x"7792",x"7793",x"7794",x"7795",x"7796",x"7797",x"7798",x"7799",x"779B",x"779C",x"779D",x"779E",x"779F",x"77A0",
x"77A1",x"77A2",x"77A4",x"77A5",x"77A6",x"77A7",x"77A8",x"77A9",x"77AA",x"77AB",x"77AC",x"77AE",x"77AF",x"77B0",x"77B1",x"77B2",
x"77B3",x"77B4",x"77B5",x"77B6",x"77B8",x"77B9",x"77BA",x"77BB",x"77BC",x"77BD",x"77BE",x"77BF",x"77C0",x"77C2",x"77C3",x"77C4",
x"77C5",x"77C6",x"77C7",x"77C8",x"77C9",x"77CA",x"77CC",x"77CD",x"77CE",x"77CF",x"77D0",x"77D1",x"77D2",x"77D3",x"77D4",x"77D6",
x"77D7",x"77D8",x"77D9",x"77DA",x"77DB",x"77DC",x"77DD",x"77DE",x"77DF",x"77E1",x"77E2",x"77E3",x"77E4",x"77E5",x"77E6",x"77E7",
x"77E8",x"77E9",x"77EA",x"77EC",x"77ED",x"77EE",x"77EF",x"77F0",x"77F1",x"77F2",x"77F3",x"77F4",x"77F5",x"77F7",x"77F8",x"77F9",
x"77FA",x"77FB",x"77FC",x"77FD",x"77FE",x"77FF",x"7800",x"7801",x"7803",x"7804",x"7805",x"7806",x"7807",x"7808",x"7809",x"780A",
x"780B",x"780C",x"780D",x"780F",x"7810",x"7811",x"7812",x"7813",x"7814",x"7815",x"7816",x"7817",x"7818",x"7819",x"781A",x"781C",
x"781D",x"781E",x"781F",x"7820",x"7821",x"7822",x"7823",x"7824",x"7825",x"7826",x"7828",x"7829",x"782A",x"782B",x"782C",x"782D",
x"782E",x"782F",x"7830",x"7831",x"7832",x"7833",x"7834",x"7836",x"7837",x"7838",x"7839",x"783A",x"783B",x"783C",x"783D",x"783E",
x"783F",x"7840",x"7841",x"7842",x"7844",x"7845",x"7846",x"7847",x"7848",x"7849",x"784A",x"784B",x"784C",x"784D",x"784E",x"784F",
x"7850",x"7852",x"7853",x"7854",x"7855",x"7856",x"7857",x"7858",x"7859",x"785A",x"785B",x"785C",x"785D",x"785E",x"785F",x"7860",
x"7862",x"7863",x"7864",x"7865",x"7866",x"7867",x"7868",x"7869",x"786A",x"786B",x"786C",x"786D",x"786E",x"786F",x"7870",x"7872",
x"7873",x"7874",x"7875",x"7876",x"7877",x"7878",x"7879",x"787A",x"787B",x"787C",x"787D",x"787E",x"787F",x"7880",x"7881",x"7883",
x"7884",x"7885",x"7886",x"7887",x"7888",x"7889",x"788A",x"788B",x"788C",x"788D",x"788E",x"788F",x"7890",x"7891",x"7892",x"7893",
x"7894",x"7896",x"7897",x"7898",x"7899",x"789A",x"789B",x"789C",x"789D",x"789E",x"789F",x"78A0",x"78A1",x"78A2",x"78A3",x"78A4",
x"78A5",x"78A6",x"78A7",x"78A8",x"78A9",x"78AB",x"78AC",x"78AD",x"78AE",x"78AF",x"78B0",x"78B1",x"78B2",x"78B3",x"78B4",x"78B5",
x"78B6",x"78B7",x"78B8",x"78B9",x"78BA",x"78BB",x"78BC",x"78BD",x"78BE",x"78BF",x"78C0",x"78C2",x"78C3",x"78C4",x"78C5",x"78C6",
x"78C7",x"78C8",x"78C9",x"78CA",x"78CB",x"78CC",x"78CD",x"78CE",x"78CF",x"78D0",x"78D1",x"78D2",x"78D3",x"78D4",x"78D5",x"78D6",
x"78D7",x"78D8",x"78D9",x"78DA",x"78DB",x"78DD",x"78DE",x"78DF",x"78E0",x"78E1",x"78E2",x"78E3",x"78E4",x"78E5",x"78E6",x"78E7",
x"78E8",x"78E9",x"78EA",x"78EB",x"78EC",x"78ED",x"78EE",x"78EF",x"78F0",x"78F1",x"78F2",x"78F3",x"78F4",x"78F5",x"78F6",x"78F7",
x"78F8",x"78F9",x"78FA",x"78FB",x"78FC",x"78FD",x"78FE",x"7900",x"7901",x"7902",x"7903",x"7904",x"7905",x"7906",x"7907",x"7908",
x"7909",x"790A",x"790B",x"790C",x"790D",x"790E",x"790F",x"7910",x"7911",x"7912",x"7913",x"7914",x"7915",x"7916",x"7917",x"7918",
x"7919",x"791A",x"791B",x"791C",x"791D",x"791E",x"791F",x"7920",x"7921",x"7922",x"7923",x"7924",x"7925",x"7926",x"7927",x"7928",
x"7929",x"792A",x"792B",x"792C",x"792D",x"792E",x"792F",x"7930",x"7931",x"7932",x"7933",x"7934",x"7935",x"7936",x"7937",x"7938",
x"7939",x"793A",x"793B",x"793C",x"793D",x"793E",x"793F",x"7940",x"7941",x"7943",x"7944",x"7945",x"7946",x"7947",x"7948",x"7949",
x"794A",x"794B",x"794C",x"794D",x"794E",x"794F",x"7950",x"7951",x"7952",x"7953",x"7954",x"7955",x"7956",x"7957",x"7958",x"7959",
x"795A",x"795B",x"795C",x"795D",x"795E",x"795F",x"7960",x"7961",x"7962",x"7963",x"7964",x"7965",x"7966",x"7967",x"7968",x"7969",
x"796A",x"796B",x"796B",x"796C",x"796D",x"796E",x"796F",x"7970",x"7971",x"7972",x"7973",x"7974",x"7975",x"7976",x"7977",x"7978",
x"7979",x"797A",x"797B",x"797C",x"797D",x"797E",x"797F",x"7980",x"7981",x"7982",x"7983",x"7984",x"7985",x"7986",x"7987",x"7988",
x"7989",x"798A",x"798B",x"798C",x"798D",x"798E",x"798F",x"7990",x"7991",x"7992",x"7993",x"7994",x"7995",x"7996",x"7997",x"7998",
x"7999",x"799A",x"799B",x"799C",x"799D",x"799E",x"799F",x"79A0",x"79A1",x"79A2",x"79A3",x"79A4",x"79A5",x"79A6",x"79A7",x"79A8",
x"79A9",x"79AA",x"79AB",x"79AC",x"79AC",x"79AD",x"79AE",x"79AF",x"79B0",x"79B1",x"79B2",x"79B3",x"79B4",x"79B5",x"79B6",x"79B7",
x"79B8",x"79B9",x"79BA",x"79BB",x"79BC",x"79BD",x"79BE",x"79BF",x"79C0",x"79C1",x"79C2",x"79C3",x"79C4",x"79C5",x"79C6",x"79C7",
x"79C8",x"79C9",x"79CA",x"79CB",x"79CC",x"79CD",x"79CD",x"79CE",x"79CF",x"79D0",x"79D1",x"79D2",x"79D3",x"79D4",x"79D5",x"79D6",
x"79D7",x"79D8",x"79D9",x"79DA",x"79DB",x"79DC",x"79DD",x"79DE",x"79DF",x"79E0",x"79E1",x"79E2",x"79E3",x"79E4",x"79E5",x"79E6",
x"79E6",x"79E7",x"79E8",x"79E9",x"79EA",x"79EB",x"79EC",x"79ED",x"79EE",x"79EF",x"79F0",x"79F1",x"79F2",x"79F3",x"79F4",x"79F5",
x"79F6",x"79F7",x"79F8",x"79F9",x"79FA",x"79FB",x"79FB",x"79FC",x"79FD",x"79FE",x"79FF",x"7A00",x"7A01",x"7A02",x"7A03",x"7A04",
x"7A05",x"7A06",x"7A07",x"7A08",x"7A09",x"7A0A",x"7A0B",x"7A0C",x"7A0D",x"7A0E",x"7A0E",x"7A0F",x"7A10",x"7A11",x"7A12",x"7A13",
x"7A14",x"7A15",x"7A16",x"7A17",x"7A18",x"7A19",x"7A1A",x"7A1B",x"7A1C",x"7A1D",x"7A1E",x"7A1E",x"7A1F",x"7A20",x"7A21",x"7A22",
x"7A23",x"7A24",x"7A25",x"7A26",x"7A27",x"7A28",x"7A29",x"7A2A",x"7A2B",x"7A2C",x"7A2D",x"7A2E",x"7A2E",x"7A2F",x"7A30",x"7A31",
x"7A32",x"7A33",x"7A34",x"7A35",x"7A36",x"7A37",x"7A38",x"7A39",x"7A3A",x"7A3B",x"7A3C",x"7A3C",x"7A3D",x"7A3E",x"7A3F",x"7A40",
x"7A41",x"7A42",x"7A43",x"7A44",x"7A45",x"7A46",x"7A47",x"7A48",x"7A49",x"7A49",x"7A4A",x"7A4B",x"7A4C",x"7A4D",x"7A4E",x"7A4F",
x"7A50",x"7A51",x"7A52",x"7A53",x"7A54",x"7A55",x"7A56",x"7A56",x"7A57",x"7A58",x"7A59",x"7A5A",x"7A5B",x"7A5C",x"7A5D",x"7A5E",
x"7A5F",x"7A60",x"7A61",x"7A61",x"7A62",x"7A63",x"7A64",x"7A65",x"7A66",x"7A67",x"7A68",x"7A69",x"7A6A",x"7A6B",x"7A6C",x"7A6D",
x"7A6D",x"7A6E",x"7A6F",x"7A70",x"7A71",x"7A72",x"7A73",x"7A74",x"7A75",x"7A76",x"7A77",x"7A78",x"7A78",x"7A79",x"7A7A",x"7A7B",
x"7A7C",x"7A7D",x"7A7E",x"7A7F",x"7A80",x"7A81",x"7A82",x"7A82",x"7A83",x"7A84",x"7A85",x"7A86",x"7A87",x"7A88",x"7A89",x"7A8A",
x"7A8B",x"7A8C",x"7A8C",x"7A8D",x"7A8E",x"7A8F",x"7A90",x"7A91",x"7A92",x"7A93",x"7A94",x"7A95",x"7A95",x"7A96",x"7A97",x"7A98",
x"7A99",x"7A9A",x"7A9B",x"7A9C",x"7A9D",x"7A9E",x"7A9F",x"7A9F",x"7AA0",x"7AA1",x"7AA2",x"7AA3",x"7AA4",x"7AA5",x"7AA6",x"7AA7",
x"7AA8",x"7AA8",x"7AA9",x"7AAA",x"7AAB",x"7AAC",x"7AAD",x"7AAE",x"7AAF",x"7AB0",x"7AB0",x"7AB1",x"7AB2",x"7AB3",x"7AB4",x"7AB5",
x"7AB6",x"7AB7",x"7AB8",x"7AB9",x"7AB9",x"7ABA",x"7ABB",x"7ABC",x"7ABD",x"7ABE",x"7ABF",x"7AC0",x"7AC1",x"7AC1",x"7AC2",x"7AC3",
x"7AC4",x"7AC5",x"7AC6",x"7AC7",x"7AC8",x"7AC9",x"7AC9",x"7ACA",x"7ACB",x"7ACC",x"7ACD",x"7ACE",x"7ACF",x"7AD0",x"7AD1",x"7AD1",
x"7AD2",x"7AD3",x"7AD4",x"7AD5",x"7AD6",x"7AD7",x"7AD8",x"7AD8",x"7AD9",x"7ADA",x"7ADB",x"7ADC",x"7ADD",x"7ADE",x"7ADF",x"7AE0",
x"7AE0",x"7AE1",x"7AE2",x"7AE3",x"7AE4",x"7AE5",x"7AE6",x"7AE7",x"7AE7",x"7AE8",x"7AE9",x"7AEA",x"7AEB",x"7AEC",x"7AED",x"7AEE",
x"7AEE",x"7AEF",x"7AF0",x"7AF1",x"7AF2",x"7AF3",x"7AF4",x"7AF5",x"7AF5",x"7AF6",x"7AF7",x"7AF8",x"7AF9",x"7AFA",x"7AFB",x"7AFC",
x"7AFC",x"7AFD",x"7AFE",x"7AFF",x"7B00",x"7B01",x"7B02",x"7B02",x"7B03",x"7B04",x"7B05",x"7B06",x"7B07",x"7B08",x"7B09",x"7B09",
x"7B0A",x"7B0B",x"7B0C",x"7B0D",x"7B0E",x"7B0F",x"7B0F",x"7B10",x"7B11",x"7B12",x"7B13",x"7B14",x"7B15",x"7B16",x"7B16",x"7B17",
x"7B18",x"7B19",x"7B1A",x"7B1B",x"7B1C",x"7B1C",x"7B1D",x"7B1E",x"7B1F",x"7B20",x"7B21",x"7B22",x"7B22",x"7B23",x"7B24",x"7B25",
x"7B26",x"7B27",x"7B28",x"7B28",x"7B29",x"7B2A",x"7B2B",x"7B2C",x"7B2D",x"7B2E",x"7B2E",x"7B2F",x"7B30",x"7B31",x"7B32",x"7B33",
x"7B33",x"7B34",x"7B35",x"7B36",x"7B37",x"7B38",x"7B39",x"7B39",x"7B3A",x"7B3B",x"7B3C",x"7B3D",x"7B3E",x"7B3F",x"7B3F",x"7B40",
x"7B41",x"7B42",x"7B43",x"7B44",x"7B44",x"7B45",x"7B46",x"7B47",x"7B48",x"7B49",x"7B4A",x"7B4A",x"7B4B",x"7B4C",x"7B4D",x"7B4E",
x"7B4F",x"7B4F",x"7B50",x"7B51",x"7B52",x"7B53",x"7B54",x"7B54",x"7B55",x"7B56",x"7B57",x"7B58",x"7B59",x"7B5A",x"7B5A",x"7B5B",
x"7B5C",x"7B5D",x"7B5E",x"7B5F",x"7B5F",x"7B60",x"7B61",x"7B62",x"7B63",x"7B64",x"7B64",x"7B65",x"7B66",x"7B67",x"7B68",x"7B69",
x"7B69",x"7B6A",x"7B6B",x"7B6C",x"7B6D",x"7B6E",x"7B6E",x"7B6F",x"7B70",x"7B71",x"7B72",x"7B73",x"7B73",x"7B74",x"7B75",x"7B76",
x"7B77",x"7B78",x"7B78",x"7B79",x"7B7A",x"7B7B",x"7B7C",x"7B7D",x"7B7D",x"7B7E",x"7B7F",x"7B80",x"7B81",x"7B81",x"7B82",x"7B83",
x"7B84",x"7B85",x"7B86",x"7B86",x"7B87",x"7B88",x"7B89",x"7B8A",x"7B8B",x"7B8B",x"7B8C",x"7B8D",x"7B8E",x"7B8F",x"7B8F",x"7B90",
x"7B91",x"7B92",x"7B93",x"7B94",x"7B94",x"7B95",x"7B96",x"7B97",x"7B98",x"7B98",x"7B99",x"7B9A",x"7B9B",x"7B9C",x"7B9D",x"7B9D",
x"7B9E",x"7B9F",x"7BA0",x"7BA1",x"7BA1",x"7BA2",x"7BA3",x"7BA4",x"7BA5",x"7BA5",x"7BA6",x"7BA7",x"7BA8",x"7BA9",x"7BAA",x"7BAA",
x"7BAB",x"7BAC",x"7BAD",x"7BAE",x"7BAE",x"7BAF",x"7BB0",x"7BB1",x"7BB2",x"7BB2",x"7BB3",x"7BB4",x"7BB5",x"7BB6",x"7BB6",x"7BB7",
x"7BB8",x"7BB9",x"7BBA",x"7BBA",x"7BBB",x"7BBC",x"7BBD",x"7BBE",x"7BBF",x"7BBF",x"7BC0",x"7BC1",x"7BC2",x"7BC3",x"7BC3",x"7BC4",
x"7BC5",x"7BC6",x"7BC7",x"7BC7",x"7BC8",x"7BC9",x"7BCA",x"7BCB",x"7BCB",x"7BCC",x"7BCD",x"7BCE",x"7BCF",x"7BCF",x"7BD0",x"7BD1",
x"7BD2",x"7BD2",x"7BD3",x"7BD4",x"7BD5",x"7BD6",x"7BD6",x"7BD7",x"7BD8",x"7BD9",x"7BDA",x"7BDA",x"7BDB",x"7BDC",x"7BDD",x"7BDE",
x"7BDE",x"7BDF",x"7BE0",x"7BE1",x"7BE2",x"7BE2",x"7BE3",x"7BE4",x"7BE5",x"7BE6",x"7BE6",x"7BE7",x"7BE8",x"7BE9",x"7BE9",x"7BEA",
x"7BEB",x"7BEC",x"7BED",x"7BED",x"7BEE",x"7BEF",x"7BF0",x"7BF1",x"7BF1",x"7BF2",x"7BF3",x"7BF4",x"7BF4",x"7BF5",x"7BF6",x"7BF7",
x"7BF8",x"7BF8",x"7BF9",x"7BFA",x"7BFB",x"7BFB",x"7BFC",x"7BFD",x"7BFE",x"7BFF",x"7BFF",x"7C00",x"7C01",x"7C02",x"7C02",x"7C03",
x"7C04",x"7C05",x"7C06",x"7C06",x"7C07",x"7C08",x"7C09",x"7C09",x"7C0A",x"7C0B",x"7C0C",x"7C0D",x"7C0D",x"7C0E",x"7C0F",x"7C10",
x"7C10",x"7C11",x"7C12",x"7C13",x"7C14",x"7C14",x"7C15",x"7C16",x"7C17",x"7C17",x"7C18",x"7C19",x"7C1A",x"7C1A",x"7C1B",x"7C1C",
x"7C1D",x"7C1E",x"7C1E",x"7C1F",x"7C20",x"7C21",x"7C21",x"7C22",x"7C23",x"7C24",x"7C24",x"7C25",x"7C26",x"7C27",x"7C27",x"7C28",
x"7C29",x"7C2A",x"7C2B",x"7C2B",x"7C2C",x"7C2D",x"7C2E",x"7C2E",x"7C2F",x"7C30",x"7C31",x"7C31",x"7C32",x"7C33",x"7C34",x"7C34",
x"7C35",x"7C36",x"7C37",x"7C37",x"7C38",x"7C39",x"7C3A",x"7C3A",x"7C3B",x"7C3C",x"7C3D",x"7C3E",x"7C3E",x"7C3F",x"7C40",x"7C41",
x"7C41",x"7C42",x"7C43",x"7C44",x"7C44",x"7C45",x"7C46",x"7C47",x"7C47",x"7C48",x"7C49",x"7C4A",x"7C4A",x"7C4B",x"7C4C",x"7C4D",
x"7C4D",x"7C4E",x"7C4F",x"7C50",x"7C50",x"7C51",x"7C52",x"7C53",x"7C53",x"7C54",x"7C55",x"7C56",x"7C56",x"7C57",x"7C58",x"7C59",
x"7C59",x"7C5A",x"7C5B",x"7C5C",x"7C5C",x"7C5D",x"7C5E",x"7C5E",x"7C5F",x"7C60",x"7C61",x"7C61",x"7C62",x"7C63",x"7C64",x"7C64",
x"7C65",x"7C66",x"7C67",x"7C67",x"7C68",x"7C69",x"7C6A",x"7C6A",x"7C6B",x"7C6C",x"7C6D",x"7C6D",x"7C6E",x"7C6F",x"7C6F",x"7C70",
x"7C71",x"7C72",x"7C72",x"7C73",x"7C74",x"7C75",x"7C75",x"7C76",x"7C77",x"7C78",x"7C78",x"7C79",x"7C7A",x"7C7A",x"7C7B",x"7C7C",
x"7C7D",x"7C7D",x"7C7E",x"7C7F",x"7C80",x"7C80",x"7C81",x"7C82",x"7C83",x"7C83",x"7C84",x"7C85",x"7C85",x"7C86",x"7C87",x"7C88",
x"7C88",x"7C89",x"7C8A",x"7C8A",x"7C8B",x"7C8C",x"7C8D",x"7C8D",x"7C8E",x"7C8F",x"7C90",x"7C90",x"7C91",x"7C92",x"7C92",x"7C93",
x"7C94",x"7C95",x"7C95",x"7C96",x"7C97",x"7C98",x"7C98",x"7C99",x"7C9A",x"7C9A",x"7C9B",x"7C9C",x"7C9D",x"7C9D",x"7C9E",x"7C9F",
x"7C9F",x"7CA0",x"7CA1",x"7CA2",x"7CA2",x"7CA3",x"7CA4",x"7CA4",x"7CA5",x"7CA6",x"7CA7",x"7CA7",x"7CA8",x"7CA9",x"7CA9",x"7CAA",
x"7CAB",x"7CAC",x"7CAC",x"7CAD",x"7CAE",x"7CAE",x"7CAF",x"7CB0",x"7CB1",x"7CB1",x"7CB2",x"7CB3",x"7CB3",x"7CB4",x"7CB5",x"7CB5",
x"7CB6",x"7CB7",x"7CB8",x"7CB8",x"7CB9",x"7CBA",x"7CBA",x"7CBB",x"7CBC",x"7CBD",x"7CBD",x"7CBE",x"7CBF",x"7CBF",x"7CC0",x"7CC1",
x"7CC1",x"7CC2",x"7CC3",x"7CC4",x"7CC4",x"7CC5",x"7CC6",x"7CC6",x"7CC7",x"7CC8",x"7CC8",x"7CC9",x"7CCA",x"7CCB",x"7CCB",x"7CCC",
x"7CCD",x"7CCD",x"7CCE",x"7CCF",x"7CCF",x"7CD0",x"7CD1",x"7CD2",x"7CD2",x"7CD3",x"7CD4",x"7CD4",x"7CD5",x"7CD6",x"7CD6",x"7CD7",
x"7CD8",x"7CD8",x"7CD9",x"7CDA",x"7CDB",x"7CDB",x"7CDC",x"7CDD",x"7CDD",x"7CDE",x"7CDF",x"7CDF",x"7CE0",x"7CE1",x"7CE1",x"7CE2",
x"7CE3",x"7CE4",x"7CE4",x"7CE5",x"7CE6",x"7CE6",x"7CE7",x"7CE8",x"7CE8",x"7CE9",x"7CEA",x"7CEA",x"7CEB",x"7CEC",x"7CEC",x"7CED",
x"7CEE",x"7CEE",x"7CEF",x"7CF0",x"7CF1",x"7CF1",x"7CF2",x"7CF3",x"7CF3",x"7CF4",x"7CF5",x"7CF5",x"7CF6",x"7CF7",x"7CF7",x"7CF8",
x"7CF9",x"7CF9",x"7CFA",x"7CFB",x"7CFB",x"7CFC",x"7CFD",x"7CFD",x"7CFE",x"7CFF",x"7CFF",x"7D00",x"7D01",x"7D02",x"7D02",x"7D03",
x"7D04",x"7D04",x"7D05",x"7D06",x"7D06",x"7D07",x"7D08",x"7D08",x"7D09",x"7D0A",x"7D0A",x"7D0B",x"7D0C",x"7D0C",x"7D0D",x"7D0E",
x"7D0E",x"7D0F",x"7D10",x"7D10",x"7D11",x"7D12",x"7D12",x"7D13",x"7D14",x"7D14",x"7D15",x"7D16",x"7D16",x"7D17",x"7D18",x"7D18",
x"7D19",x"7D1A",x"7D1A",x"7D1B",x"7D1C",x"7D1C",x"7D1D",x"7D1E",x"7D1E",x"7D1F",x"7D20",x"7D20",x"7D21",x"7D22",x"7D22",x"7D23",
x"7D24",x"7D24",x"7D25",x"7D26",x"7D26",x"7D27",x"7D28",x"7D28",x"7D29",x"7D29",x"7D2A",x"7D2B",x"7D2B",x"7D2C",x"7D2D",x"7D2D",
x"7D2E",x"7D2F",x"7D2F",x"7D30",x"7D31",x"7D31",x"7D32",x"7D33",x"7D33",x"7D34",x"7D35",x"7D35",x"7D36",x"7D37",x"7D37",x"7D38",
x"7D39",x"7D39",x"7D3A",x"7D3A",x"7D3B",x"7D3C",x"7D3C",x"7D3D",x"7D3E",x"7D3E",x"7D3F",x"7D40",x"7D40",x"7D41",x"7D42",x"7D42",
x"7D43",x"7D44",x"7D44",x"7D45",x"7D45",x"7D46",x"7D47",x"7D47",x"7D48",x"7D49",x"7D49",x"7D4A",x"7D4B",x"7D4B",x"7D4C",x"7D4D",
x"7D4D",x"7D4E",x"7D4E",x"7D4F",x"7D50",x"7D50",x"7D51",x"7D52",x"7D52",x"7D53",x"7D54",x"7D54",x"7D55",x"7D56",x"7D56",x"7D57",
x"7D57",x"7D58",x"7D59",x"7D59",x"7D5A",x"7D5B",x"7D5B",x"7D5C",x"7D5C",x"7D5D",x"7D5E",x"7D5E",x"7D5F",x"7D60",x"7D60",x"7D61",
x"7D62",x"7D62",x"7D63",x"7D63",x"7D64",x"7D65",x"7D65",x"7D66",x"7D67",x"7D67",x"7D68",x"7D68",x"7D69",x"7D6A",x"7D6A",x"7D6B",
x"7D6C",x"7D6C",x"7D6D",x"7D6E",x"7D6E",x"7D6F",x"7D6F",x"7D70",x"7D71",x"7D71",x"7D72",x"7D73",x"7D73",x"7D74",x"7D74",x"7D75",
x"7D76",x"7D76",x"7D77",x"7D77",x"7D78",x"7D79",x"7D79",x"7D7A",x"7D7B",x"7D7B",x"7D7C",x"7D7C",x"7D7D",x"7D7E",x"7D7E",x"7D7F",
x"7D80",x"7D80",x"7D81",x"7D81",x"7D82",x"7D83",x"7D83",x"7D84",x"7D84",x"7D85",x"7D86",x"7D86",x"7D87",x"7D88",x"7D88",x"7D89",
x"7D89",x"7D8A",x"7D8B",x"7D8B",x"7D8C",x"7D8C",x"7D8D",x"7D8E",x"7D8E",x"7D8F",x"7D90",x"7D90",x"7D91",x"7D91",x"7D92",x"7D93",
x"7D93",x"7D94",x"7D94",x"7D95",x"7D96",x"7D96",x"7D97",x"7D97",x"7D98",x"7D99",x"7D99",x"7D9A",x"7D9A",x"7D9B",x"7D9C",x"7D9C",
x"7D9D",x"7D9D",x"7D9E",x"7D9F",x"7D9F",x"7DA0",x"7DA0",x"7DA1",x"7DA2",x"7DA2",x"7DA3",x"7DA3",x"7DA4",x"7DA5",x"7DA5",x"7DA6",
x"7DA6",x"7DA7",x"7DA8",x"7DA8",x"7DA9",x"7DA9",x"7DAA",x"7DAB",x"7DAB",x"7DAC",x"7DAC",x"7DAD",x"7DAE",x"7DAE",x"7DAF",x"7DAF",
x"7DB0",x"7DB1",x"7DB1",x"7DB2",x"7DB2",x"7DB3",x"7DB4",x"7DB4",x"7DB5",x"7DB5",x"7DB6",x"7DB7",x"7DB7",x"7DB8",x"7DB8",x"7DB9",
x"7DB9",x"7DBA",x"7DBB",x"7DBB",x"7DBC",x"7DBC",x"7DBD",x"7DBE",x"7DBE",x"7DBF",x"7DBF",x"7DC0",x"7DC1",x"7DC1",x"7DC2",x"7DC2",
x"7DC3",x"7DC3",x"7DC4",x"7DC5",x"7DC5",x"7DC6",x"7DC6",x"7DC7",x"7DC8",x"7DC8",x"7DC9",x"7DC9",x"7DCA",x"7DCA",x"7DCB",x"7DCC",
x"7DCC",x"7DCD",x"7DCD",x"7DCE",x"7DCE",x"7DCF",x"7DD0",x"7DD0",x"7DD1",x"7DD1",x"7DD2",x"7DD3",x"7DD3",x"7DD4",x"7DD4",x"7DD5",
x"7DD5",x"7DD6",x"7DD7",x"7DD7",x"7DD8",x"7DD8",x"7DD9",x"7DD9",x"7DDA",x"7DDB",x"7DDB",x"7DDC",x"7DDC",x"7DDD",x"7DDD",x"7DDE",
x"7DDF",x"7DDF",x"7DE0",x"7DE0",x"7DE1",x"7DE1",x"7DE2",x"7DE3",x"7DE3",x"7DE4",x"7DE4",x"7DE5",x"7DE5",x"7DE6",x"7DE7",x"7DE7",
x"7DE8",x"7DE8",x"7DE9",x"7DE9",x"7DEA",x"7DEA",x"7DEB",x"7DEC",x"7DEC",x"7DED",x"7DED",x"7DEE",x"7DEE",x"7DEF",x"7DF0",x"7DF0",
x"7DF1",x"7DF1",x"7DF2",x"7DF2",x"7DF3",x"7DF3",x"7DF4",x"7DF5",x"7DF5",x"7DF6",x"7DF6",x"7DF7",x"7DF7",x"7DF8",x"7DF8",x"7DF9",
x"7DFA",x"7DFA",x"7DFB",x"7DFB",x"7DFC",x"7DFC",x"7DFD",x"7DFD",x"7DFE",x"7DFF",x"7DFF",x"7E00",x"7E00",x"7E01",x"7E01",x"7E02",
x"7E02",x"7E03",x"7E04",x"7E04",x"7E05",x"7E05",x"7E06",x"7E06",x"7E07",x"7E07",x"7E08",x"7E09",x"7E09",x"7E0A",x"7E0A",x"7E0B",
x"7E0B",x"7E0C",x"7E0C",x"7E0D",x"7E0D",x"7E0E",x"7E0F",x"7E0F",x"7E10",x"7E10",x"7E11",x"7E11",x"7E12",x"7E12",x"7E13",x"7E13",
x"7E14",x"7E15",x"7E15",x"7E16",x"7E16",x"7E17",x"7E17",x"7E18",x"7E18",x"7E19",x"7E19",x"7E1A",x"7E1A",x"7E1B",x"7E1C",x"7E1C",
x"7E1D",x"7E1D",x"7E1E",x"7E1E",x"7E1F",x"7E1F",x"7E20",x"7E20",x"7E21",x"7E21",x"7E22",x"7E22",x"7E23",x"7E24",x"7E24",x"7E25",
x"7E25",x"7E26",x"7E26",x"7E27",x"7E27",x"7E28",x"7E28",x"7E29",x"7E29",x"7E2A",x"7E2A",x"7E2B",x"7E2C",x"7E2C",x"7E2D",x"7E2D",
x"7E2E",x"7E2E",x"7E2F",x"7E2F",x"7E30",x"7E30",x"7E31",x"7E31",x"7E32",x"7E32",x"7E33",x"7E33",x"7E34",x"7E34",x"7E35",x"7E36",
x"7E36",x"7E37",x"7E37",x"7E38",x"7E38",x"7E39",x"7E39",x"7E3A",x"7E3A",x"7E3B",x"7E3B",x"7E3C",x"7E3C",x"7E3D",x"7E3D",x"7E3E",
x"7E3E",x"7E3F",x"7E3F",x"7E40",x"7E40",x"7E41",x"7E41",x"7E42",x"7E42",x"7E43",x"7E44",x"7E44",x"7E45",x"7E45",x"7E46",x"7E46",
x"7E47",x"7E47",x"7E48",x"7E48",x"7E49",x"7E49",x"7E4A",x"7E4A",x"7E4B",x"7E4B",x"7E4C",x"7E4C",x"7E4D",x"7E4D",x"7E4E",x"7E4E",
x"7E4F",x"7E4F",x"7E50",x"7E50",x"7E51",x"7E51",x"7E52",x"7E52",x"7E53",x"7E53",x"7E54",x"7E54",x"7E55",x"7E55",x"7E56",x"7E56",
x"7E57",x"7E57",x"7E58",x"7E58",x"7E59",x"7E59",x"7E5A",x"7E5A",x"7E5B",x"7E5B",x"7E5C",x"7E5C",x"7E5D",x"7E5D",x"7E5E",x"7E5E",
x"7E5F",x"7E5F",x"7E60",x"7E60",x"7E61",x"7E61",x"7E62",x"7E62",x"7E63",x"7E63",x"7E64",x"7E64",x"7E65",x"7E65",x"7E66",x"7E66",
x"7E67",x"7E67",x"7E68",x"7E68",x"7E69",x"7E69",x"7E6A",x"7E6A",x"7E6B",x"7E6B",x"7E6C",x"7E6C",x"7E6D",x"7E6D",x"7E6E",x"7E6E",
x"7E6F",x"7E6F",x"7E70",x"7E70",x"7E71",x"7E71",x"7E72",x"7E72",x"7E73",x"7E73",x"7E74",x"7E74",x"7E75",x"7E75",x"7E76",x"7E76",
x"7E77",x"7E77",x"7E77",x"7E78",x"7E78",x"7E79",x"7E79",x"7E7A",x"7E7A",x"7E7B",x"7E7B",x"7E7C",x"7E7C",x"7E7D",x"7E7D",x"7E7E",
x"7E7E",x"7E7F",x"7E7F",x"7E80",x"7E80",x"7E81",x"7E81",x"7E82",x"7E82",x"7E83",x"7E83",x"7E83",x"7E84",x"7E84",x"7E85",x"7E85",
x"7E86",x"7E86",x"7E87",x"7E87",x"7E88",x"7E88",x"7E89",x"7E89",x"7E8A",x"7E8A",x"7E8B",x"7E8B",x"7E8C",x"7E8C",x"7E8D",x"7E8D",
x"7E8D",x"7E8E",x"7E8E",x"7E8F",x"7E8F",x"7E90",x"7E90",x"7E91",x"7E91",x"7E92",x"7E92",x"7E93",x"7E93",x"7E94",x"7E94",x"7E94",
x"7E95",x"7E95",x"7E96",x"7E96",x"7E97",x"7E97",x"7E98",x"7E98",x"7E99",x"7E99",x"7E9A",x"7E9A",x"7E9B",x"7E9B",x"7E9B",x"7E9C",
x"7E9C",x"7E9D",x"7E9D",x"7E9E",x"7E9E",x"7E9F",x"7E9F",x"7EA0",x"7EA0",x"7EA0",x"7EA1",x"7EA1",x"7EA2",x"7EA2",x"7EA3",x"7EA3",
x"7EA4",x"7EA4",x"7EA5",x"7EA5",x"7EA6",x"7EA6",x"7EA6",x"7EA7",x"7EA7",x"7EA8",x"7EA8",x"7EA9",x"7EA9",x"7EAA",x"7EAA",x"7EAA",
x"7EAB",x"7EAB",x"7EAC",x"7EAC",x"7EAD",x"7EAD",x"7EAE",x"7EAE",x"7EAF",x"7EAF",x"7EAF",x"7EB0",x"7EB0",x"7EB1",x"7EB1",x"7EB2",
x"7EB2",x"7EB3",x"7EB3",x"7EB3",x"7EB4",x"7EB4",x"7EB5",x"7EB5",x"7EB6",x"7EB6",x"7EB7",x"7EB7",x"7EB7",x"7EB8",x"7EB8",x"7EB9",
x"7EB9",x"7EBA",x"7EBA",x"7EBB",x"7EBB",x"7EBB",x"7EBC",x"7EBC",x"7EBD",x"7EBD",x"7EBE",x"7EBE",x"7EBF",x"7EBF",x"7EBF",x"7EC0",
x"7EC0",x"7EC1",x"7EC1",x"7EC2",x"7EC2",x"7EC2",x"7EC3",x"7EC3",x"7EC4",x"7EC4",x"7EC5",x"7EC5",x"7EC5",x"7EC6",x"7EC6",x"7EC7",
x"7EC7",x"7EC8",x"7EC8",x"7EC9",x"7EC9",x"7EC9",x"7ECA",x"7ECA",x"7ECB",x"7ECB",x"7ECC",x"7ECC",x"7ECC",x"7ECD",x"7ECD",x"7ECE",
x"7ECE",x"7ECF",x"7ECF",x"7ECF",x"7ED0",x"7ED0",x"7ED1",x"7ED1",x"7ED2",x"7ED2",x"7ED2",x"7ED3",x"7ED3",x"7ED4",x"7ED4",x"7ED4",
x"7ED5",x"7ED5",x"7ED6",x"7ED6",x"7ED7",x"7ED7",x"7ED7",x"7ED8",x"7ED8",x"7ED9",x"7ED9",x"7EDA",x"7EDA",x"7EDA",x"7EDB",x"7EDB",
x"7EDC",x"7EDC",x"7EDC",x"7EDD",x"7EDD",x"7EDE",x"7EDE",x"7EDF",x"7EDF",x"7EDF",x"7EE0",x"7EE0",x"7EE1",x"7EE1",x"7EE1",x"7EE2",
x"7EE2",x"7EE3",x"7EE3",x"7EE4",x"7EE4",x"7EE4",x"7EE5",x"7EE5",x"7EE6",x"7EE6",x"7EE6",x"7EE7",x"7EE7",x"7EE8",x"7EE8",x"7EE8",
x"7EE9",x"7EE9",x"7EEA",x"7EEA",x"7EEA",x"7EEB",x"7EEB",x"7EEC",x"7EEC",x"7EED",x"7EED",x"7EED",x"7EEE",x"7EEE",x"7EEF",x"7EEF",
x"7EEF",x"7EF0",x"7EF0",x"7EF1",x"7EF1",x"7EF1",x"7EF2",x"7EF2",x"7EF3",x"7EF3",x"7EF3",x"7EF4",x"7EF4",x"7EF5",x"7EF5",x"7EF5",
x"7EF6",x"7EF6",x"7EF7",x"7EF7",x"7EF7",x"7EF8",x"7EF8",x"7EF9",x"7EF9",x"7EF9",x"7EFA",x"7EFA",x"7EFB",x"7EFB",x"7EFB",x"7EFC",
x"7EFC",x"7EFD",x"7EFD",x"7EFD",x"7EFE",x"7EFE",x"7EFE",x"7EFF",x"7EFF",x"7F00",x"7F00",x"7F00",x"7F01",x"7F01",x"7F02",x"7F02",
x"7F02",x"7F03",x"7F03",x"7F04",x"7F04",x"7F04",x"7F05",x"7F05",x"7F05",x"7F06",x"7F06",x"7F07",x"7F07",x"7F07",x"7F08",x"7F08",
x"7F09",x"7F09",x"7F09",x"7F0A",x"7F0A",x"7F0A",x"7F0B",x"7F0B",x"7F0C",x"7F0C",x"7F0C",x"7F0D",x"7F0D",x"7F0E",x"7F0E",x"7F0E",
x"7F0F",x"7F0F",x"7F0F",x"7F10",x"7F10",x"7F11",x"7F11",x"7F11",x"7F12",x"7F12",x"7F12",x"7F13",x"7F13",x"7F14",x"7F14",x"7F14",
x"7F15",x"7F15",x"7F15",x"7F16",x"7F16",x"7F17",x"7F17",x"7F17",x"7F18",x"7F18",x"7F18",x"7F19",x"7F19",x"7F1A",x"7F1A",x"7F1A",
x"7F1B",x"7F1B",x"7F1B",x"7F1C",x"7F1C",x"7F1D",x"7F1D",x"7F1D",x"7F1E",x"7F1E",x"7F1E",x"7F1F",x"7F1F",x"7F1F",x"7F20",x"7F20",
x"7F21",x"7F21",x"7F21",x"7F22",x"7F22",x"7F22",x"7F23",x"7F23",x"7F23",x"7F24",x"7F24",x"7F25",x"7F25",x"7F25",x"7F26",x"7F26",
x"7F26",x"7F27",x"7F27",x"7F27",x"7F28",x"7F28",x"7F29",x"7F29",x"7F29",x"7F2A",x"7F2A",x"7F2A",x"7F2B",x"7F2B",x"7F2B",x"7F2C",
x"7F2C",x"7F2C",x"7F2D",x"7F2D",x"7F2E",x"7F2E",x"7F2E",x"7F2F",x"7F2F",x"7F2F",x"7F30",x"7F30",x"7F30",x"7F31",x"7F31",x"7F31",
x"7F32",x"7F32",x"7F32",x"7F33",x"7F33",x"7F34",x"7F34",x"7F34",x"7F35",x"7F35",x"7F35",x"7F36",x"7F36",x"7F36",x"7F37",x"7F37",
x"7F37",x"7F38",x"7F38",x"7F38",x"7F39",x"7F39",x"7F39",x"7F3A",x"7F3A",x"7F3A",x"7F3B",x"7F3B",x"7F3B",x"7F3C",x"7F3C",x"7F3D",
x"7F3D",x"7F3D",x"7F3E",x"7F3E",x"7F3E",x"7F3F",x"7F3F",x"7F3F",x"7F40",x"7F40",x"7F40",x"7F41",x"7F41",x"7F41",x"7F42",x"7F42",
x"7F42",x"7F43",x"7F43",x"7F43",x"7F44",x"7F44",x"7F44",x"7F45",x"7F45",x"7F45",x"7F46",x"7F46",x"7F46",x"7F47",x"7F47",x"7F47",
x"7F48",x"7F48",x"7F48",x"7F49",x"7F49",x"7F49",x"7F4A",x"7F4A",x"7F4A",x"7F4B",x"7F4B",x"7F4B",x"7F4C",x"7F4C",x"7F4C",x"7F4D",
x"7F4D",x"7F4D",x"7F4E",x"7F4E",x"7F4E",x"7F4F",x"7F4F",x"7F4F",x"7F50",x"7F50",x"7F50",x"7F50",x"7F51",x"7F51",x"7F51",x"7F52",
x"7F52",x"7F52",x"7F53",x"7F53",x"7F53",x"7F54",x"7F54",x"7F54",x"7F55",x"7F55",x"7F55",x"7F56",x"7F56",x"7F56",x"7F57",x"7F57",
x"7F57",x"7F58",x"7F58",x"7F58",x"7F58",x"7F59",x"7F59",x"7F59",x"7F5A",x"7F5A",x"7F5A",x"7F5B",x"7F5B",x"7F5B",x"7F5C",x"7F5C",
x"7F5C",x"7F5D",x"7F5D",x"7F5D",x"7F5E",x"7F5E",x"7F5E",x"7F5E",x"7F5F",x"7F5F",x"7F5F",x"7F60",x"7F60",x"7F60",x"7F61",x"7F61",
x"7F61",x"7F62",x"7F62",x"7F62",x"7F62",x"7F63",x"7F63",x"7F63",x"7F64",x"7F64",x"7F64",x"7F65",x"7F65",x"7F65",x"7F65",x"7F66",
x"7F66",x"7F66",x"7F67",x"7F67",x"7F67",x"7F68",x"7F68",x"7F68",x"7F69",x"7F69",x"7F69",x"7F69",x"7F6A",x"7F6A",x"7F6A",x"7F6B",
x"7F6B",x"7F6B",x"7F6C",x"7F6C",x"7F6C",x"7F6C",x"7F6D",x"7F6D",x"7F6D",x"7F6E",x"7F6E",x"7F6E",x"7F6E",x"7F6F",x"7F6F",x"7F6F",
x"7F70",x"7F70",x"7F70",x"7F71",x"7F71",x"7F71",x"7F71",x"7F72",x"7F72",x"7F72",x"7F73",x"7F73",x"7F73",x"7F73",x"7F74",x"7F74",
x"7F74",x"7F75",x"7F75",x"7F75",x"7F75",x"7F76",x"7F76",x"7F76",x"7F77",x"7F77",x"7F77",x"7F77",x"7F78",x"7F78",x"7F78",x"7F79",
x"7F79",x"7F79",x"7F79",x"7F7A",x"7F7A",x"7F7A",x"7F7B",x"7F7B",x"7F7B",x"7F7B",x"7F7C",x"7F7C",x"7F7C",x"7F7D",x"7F7D",x"7F7D",
x"7F7D",x"7F7E",x"7F7E",x"7F7E",x"7F7F",x"7F7F",x"7F7F",x"7F7F",x"7F80",x"7F80",x"7F80",x"7F80",x"7F81",x"7F81",x"7F81",x"7F82",
x"7F82",x"7F82",x"7F82",x"7F83",x"7F83",x"7F83",x"7F83",x"7F84",x"7F84",x"7F84",x"7F85",x"7F85",x"7F85",x"7F85",x"7F86",x"7F86",
x"7F86",x"7F86",x"7F87",x"7F87",x"7F87",x"7F88",x"7F88",x"7F88",x"7F88",x"7F89",x"7F89",x"7F89",x"7F89",x"7F8A",x"7F8A",x"7F8A",
x"7F8A",x"7F8B",x"7F8B",x"7F8B",x"7F8C",x"7F8C",x"7F8C",x"7F8C",x"7F8D",x"7F8D",x"7F8D",x"7F8D",x"7F8E",x"7F8E",x"7F8E",x"7F8E",
x"7F8F",x"7F8F",x"7F8F",x"7F8F",x"7F90",x"7F90",x"7F90",x"7F90",x"7F91",x"7F91",x"7F91",x"7F91",x"7F92",x"7F92",x"7F92",x"7F93",
x"7F93",x"7F93",x"7F93",x"7F94",x"7F94",x"7F94",x"7F94",x"7F95",x"7F95",x"7F95",x"7F95",x"7F96",x"7F96",x"7F96",x"7F96",x"7F97",
x"7F97",x"7F97",x"7F97",x"7F98",x"7F98",x"7F98",x"7F98",x"7F99",x"7F99",x"7F99",x"7F99",x"7F9A",x"7F9A",x"7F9A",x"7F9A",x"7F9B",
x"7F9B",x"7F9B",x"7F9B",x"7F9C",x"7F9C",x"7F9C",x"7F9C",x"7F9C",x"7F9D",x"7F9D",x"7F9D",x"7F9D",x"7F9E",x"7F9E",x"7F9E",x"7F9E",
x"7F9F",x"7F9F",x"7F9F",x"7F9F",x"7FA0",x"7FA0",x"7FA0",x"7FA0",x"7FA1",x"7FA1",x"7FA1",x"7FA1",x"7FA2",x"7FA2",x"7FA2",x"7FA2",
x"7FA2",x"7FA3",x"7FA3",x"7FA3",x"7FA3",x"7FA4",x"7FA4",x"7FA4",x"7FA4",x"7FA5",x"7FA5",x"7FA5",x"7FA5",x"7FA6",x"7FA6",x"7FA6",
x"7FA6",x"7FA6",x"7FA7",x"7FA7",x"7FA7",x"7FA7",x"7FA8",x"7FA8",x"7FA8",x"7FA8",x"7FA9",x"7FA9",x"7FA9",x"7FA9",x"7FA9",x"7FAA",
x"7FAA",x"7FAA",x"7FAA",x"7FAB",x"7FAB",x"7FAB",x"7FAB",x"7FAB",x"7FAC",x"7FAC",x"7FAC",x"7FAC",x"7FAD",x"7FAD",x"7FAD",x"7FAD",
x"7FAD",x"7FAE",x"7FAE",x"7FAE",x"7FAE",x"7FAF",x"7FAF",x"7FAF",x"7FAF",x"7FAF",x"7FB0",x"7FB0",x"7FB0",x"7FB0",x"7FB1",x"7FB1",
x"7FB1",x"7FB1",x"7FB1",x"7FB2",x"7FB2",x"7FB2",x"7FB2",x"7FB2",x"7FB3",x"7FB3",x"7FB3",x"7FB3",x"7FB4",x"7FB4",x"7FB4",x"7FB4",
x"7FB4",x"7FB5",x"7FB5",x"7FB5",x"7FB5",x"7FB5",x"7FB6",x"7FB6",x"7FB6",x"7FB6",x"7FB6",x"7FB7",x"7FB7",x"7FB7",x"7FB7",x"7FB8",
x"7FB8",x"7FB8",x"7FB8",x"7FB8",x"7FB9",x"7FB9",x"7FB9",x"7FB9",x"7FB9",x"7FBA",x"7FBA",x"7FBA",x"7FBA",x"7FBA",x"7FBB",x"7FBB",
x"7FBB",x"7FBB",x"7FBB",x"7FBC",x"7FBC",x"7FBC",x"7FBC",x"7FBC",x"7FBD",x"7FBD",x"7FBD",x"7FBD",x"7FBD",x"7FBE",x"7FBE",x"7FBE",
x"7FBE",x"7FBE",x"7FBF",x"7FBF",x"7FBF",x"7FBF",x"7FBF",x"7FC0",x"7FC0",x"7FC0",x"7FC0",x"7FC0",x"7FC1",x"7FC1",x"7FC1",x"7FC1",
x"7FC1",x"7FC2",x"7FC2",x"7FC2",x"7FC2",x"7FC2",x"7FC2",x"7FC3",x"7FC3",x"7FC3",x"7FC3",x"7FC3",x"7FC4",x"7FC4",x"7FC4",x"7FC4",
x"7FC4",x"7FC5",x"7FC5",x"7FC5",x"7FC5",x"7FC5",x"7FC6",x"7FC6",x"7FC6",x"7FC6",x"7FC6",x"7FC6",x"7FC7",x"7FC7",x"7FC7",x"7FC7",
x"7FC7",x"7FC8",x"7FC8",x"7FC8",x"7FC8",x"7FC8",x"7FC8",x"7FC9",x"7FC9",x"7FC9",x"7FC9",x"7FC9",x"7FCA",x"7FCA",x"7FCA",x"7FCA",
x"7FCA",x"7FCA",x"7FCB",x"7FCB",x"7FCB",x"7FCB",x"7FCB",x"7FCB",x"7FCC",x"7FCC",x"7FCC",x"7FCC",x"7FCC",x"7FCD",x"7FCD",x"7FCD",
x"7FCD",x"7FCD",x"7FCD",x"7FCE",x"7FCE",x"7FCE",x"7FCE",x"7FCE",x"7FCE",x"7FCF",x"7FCF",x"7FCF",x"7FCF",x"7FCF",x"7FCF",x"7FD0",
x"7FD0",x"7FD0",x"7FD0",x"7FD0",x"7FD0",x"7FD1",x"7FD1",x"7FD1",x"7FD1",x"7FD1",x"7FD1",x"7FD2",x"7FD2",x"7FD2",x"7FD2",x"7FD2",
x"7FD2",x"7FD3",x"7FD3",x"7FD3",x"7FD3",x"7FD3",x"7FD3",x"7FD4",x"7FD4",x"7FD4",x"7FD4",x"7FD4",x"7FD4",x"7FD5",x"7FD5",x"7FD5",
x"7FD5",x"7FD5",x"7FD5",x"7FD6",x"7FD6",x"7FD6",x"7FD6",x"7FD6",x"7FD6",x"7FD6",x"7FD7",x"7FD7",x"7FD7",x"7FD7",x"7FD7",x"7FD7",
x"7FD8",x"7FD8",x"7FD8",x"7FD8",x"7FD8",x"7FD8",x"7FD8",x"7FD9",x"7FD9",x"7FD9",x"7FD9",x"7FD9",x"7FD9",x"7FDA",x"7FDA",x"7FDA",
x"7FDA",x"7FDA",x"7FDA",x"7FDA",x"7FDB",x"7FDB",x"7FDB",x"7FDB",x"7FDB",x"7FDB",x"7FDB",x"7FDC",x"7FDC",x"7FDC",x"7FDC",x"7FDC",
x"7FDC",x"7FDC",x"7FDD",x"7FDD",x"7FDD",x"7FDD",x"7FDD",x"7FDD",x"7FDD",x"7FDE",x"7FDE",x"7FDE",x"7FDE",x"7FDE",x"7FDE",x"7FDE",
x"7FDF",x"7FDF",x"7FDF",x"7FDF",x"7FDF",x"7FDF",x"7FDF",x"7FE0",x"7FE0",x"7FE0",x"7FE0",x"7FE0",x"7FE0",x"7FE0",x"7FE1",x"7FE1",
x"7FE1",x"7FE1",x"7FE1",x"7FE1",x"7FE1",x"7FE1",x"7FE2",x"7FE2",x"7FE2",x"7FE2",x"7FE2",x"7FE2",x"7FE2",x"7FE3",x"7FE3",x"7FE3",
x"7FE3",x"7FE3",x"7FE3",x"7FE3",x"7FE3",x"7FE4",x"7FE4",x"7FE4",x"7FE4",x"7FE4",x"7FE4",x"7FE4",x"7FE4",x"7FE5",x"7FE5",x"7FE5",
x"7FE5",x"7FE5",x"7FE5",x"7FE5",x"7FE5",x"7FE6",x"7FE6",x"7FE6",x"7FE6",x"7FE6",x"7FE6",x"7FE6",x"7FE6",x"7FE7",x"7FE7",x"7FE7",
x"7FE7",x"7FE7",x"7FE7",x"7FE7",x"7FE7",x"7FE8",x"7FE8",x"7FE8",x"7FE8",x"7FE8",x"7FE8",x"7FE8",x"7FE8",x"7FE8",x"7FE9",x"7FE9",
x"7FE9",x"7FE9",x"7FE9",x"7FE9",x"7FE9",x"7FE9",x"7FE9",x"7FEA",x"7FEA",x"7FEA",x"7FEA",x"7FEA",x"7FEA",x"7FEA",x"7FEA",x"7FEA",
x"7FEB",x"7FEB",x"7FEB",x"7FEB",x"7FEB",x"7FEB",x"7FEB",x"7FEB",x"7FEB",x"7FEC",x"7FEC",x"7FEC",x"7FEC",x"7FEC",x"7FEC",x"7FEC",
x"7FEC",x"7FEC",x"7FED",x"7FED",x"7FED",x"7FED",x"7FED",x"7FED",x"7FED",x"7FED",x"7FED",x"7FED",x"7FEE",x"7FEE",x"7FEE",x"7FEE",
x"7FEE",x"7FEE",x"7FEE",x"7FEE",x"7FEE",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",x"7FEF",
x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF0",x"7FF1",x"7FF1",x"7FF1",x"7FF1",x"7FF1",x"7FF1",
x"7FF1",x"7FF1",x"7FF1",x"7FF1",x"7FF1",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",x"7FF2",
x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF3",x"7FF4",x"7FF4",x"7FF4",x"7FF4",
x"7FF4",x"7FF4",x"7FF4",x"7FF4",x"7FF4",x"7FF4",x"7FF4",x"7FF4",x"7FF5",x"7FF5",x"7FF5",x"7FF5",x"7FF5",x"7FF5",x"7FF5",x"7FF5",
x"7FF5",x"7FF5",x"7FF5",x"7FF5",x"7FF5",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",x"7FF6",
x"7FF6",x"7FF6",x"7FF6",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",x"7FF7",
x"7FF7",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",x"7FF8",
x"7FF8",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",x"7FF9",
x"7FF9",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFA",
x"7FFA",x"7FFA",x"7FFA",x"7FFA",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",
x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFB",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",
x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",x"7FFC",
x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",
x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFD",x"7FFE",x"7FFE",x"7FFE",
x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",
x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",
x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFE",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",
x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",
x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",
x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF",x"7FFF" );
       
-- Vivado specific attributes to force use of BlockRAM   
attribute rom_style : string;
attribute rom_style of rom : signal is "block";
   
    
begin

  process (CLK)
  begin
    if (CLK'event and CLK = '1') then
      dataA <= rom(to_integer(unsigned(ADDRESS_A)));
    end if;
  end process;
  
  process (CLK)
  begin
    if (CLK'event and CLK = '1') then
      DATAOUT_A <= dataA;
    end if;
  end process;
  
  

  process (CLK)
  begin
    if (CLK'event and CLK = '1') then
      dataB <= rom(to_integer(unsigned(ADDRESS_B)));
    end if;
  end process;
  
  process (CLK)
  begin
    if (CLK'event and CLK = '1') then
      DATAOUT_B <= dataB;
    end if;
  end process;
  


end architecture arcdpROM;
-----------------------------------------------------------------
--   End of File: dpROM16_v1_0.vhd
-----------------------------------------------------------------


